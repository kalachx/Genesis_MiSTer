`timescale 1ns / 1ps


/* This file is part of JT12 modification adding high precission audio
   mode called FM Overdrive
 
    JT12 program is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.

    JT12 program is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.

    You should have received a copy of the GNU General Public License
    along with JT12.  If not, see <http://www.gnu.org/licenses/>.

    Based on Sauraen VHDL version of OPN/OPN2, which is based on die shots.

    Author: Jose Tejada Gomez. Twitter: @topapate
    Version: 1.0
    Date: 27-1-2017 

*/

// altera message_off 10030

module jt12_exprom_hd
(
    input [19:0] addr,
    input clk, 
    input clk_en,
    input fmo_exprom,
    output reg [21:0] exp
);

always @ (posedge clk) if(clk_en)
    case (fmo_exprom)
        1'b0: // exponent
            case (addr[19:8])
                12'd0000: exp <= 22'd4192885;
                12'd0001: exp <= 22'd4191465;
                12'd0002: exp <= 22'd4190046;
                12'd0003: exp <= 22'd4188628;
                12'd0004: exp <= 22'd4187209;
                12'd0005: exp <= 22'd4185791;
                12'd0006: exp <= 22'd4184373;
                12'd0007: exp <= 22'd4182955;
                12'd0008: exp <= 22'd4181538;
                12'd0009: exp <= 22'd4180120;
                12'd0010: exp <= 22'd4178703;
                12'd0011: exp <= 22'd4177286;
                12'd0012: exp <= 22'd4175870;
                12'd0013: exp <= 22'd4174454;
                12'd0014: exp <= 22'd4173038;
                12'd0015: exp <= 22'd4171622;
                12'd0016: exp <= 22'd4170206;
                12'd0017: exp <= 22'd4168791;
                12'd0018: exp <= 22'd4167376;
                12'd0019: exp <= 22'd4165961;
                12'd0020: exp <= 22'd4164546;
                12'd0021: exp <= 22'd4163132;
                12'd0022: exp <= 22'd4161717;
                12'd0023: exp <= 22'd4160304;
                12'd0024: exp <= 22'd4158890;
                12'd0025: exp <= 22'd4157476;
                12'd0026: exp <= 22'd4156063;
                12'd0027: exp <= 22'd4154650;
                12'd0028: exp <= 22'd4153237;
                12'd0029: exp <= 22'd4151825;
                12'd0030: exp <= 22'd4150413;
                12'd0031: exp <= 22'd4149001;
                12'd0032: exp <= 22'd4147589;
                12'd0033: exp <= 22'd4146177;
                12'd0034: exp <= 22'd4144766;
                12'd0035: exp <= 22'd4143355;
                12'd0036: exp <= 22'd4141944;
                12'd0037: exp <= 22'd4140534;
                12'd0038: exp <= 22'd4139123;
                12'd0039: exp <= 22'd4137713;
                12'd0040: exp <= 22'd4136303;
                12'd0041: exp <= 22'd4134894;
                12'd0042: exp <= 22'd4133484;
                12'd0043: exp <= 22'd4132075;
                12'd0044: exp <= 22'd4130666;
                12'd0045: exp <= 22'd4129257;
                12'd0046: exp <= 22'd4127849;
                12'd0047: exp <= 22'd4126441;
                12'd0048: exp <= 22'd4125033;
                12'd0049: exp <= 22'd4123625;
                12'd0050: exp <= 22'd4122218;
                12'd0051: exp <= 22'd4120810;
                12'd0052: exp <= 22'd4119403;
                12'd0053: exp <= 22'd4117997;
                12'd0054: exp <= 22'd4116590;
                12'd0055: exp <= 22'd4115184;
                12'd0056: exp <= 22'd4113778;
                12'd0057: exp <= 22'd4112372;
                12'd0058: exp <= 22'd4110966;
                12'd0059: exp <= 22'd4109561;
                12'd0060: exp <= 22'd4108156;
                12'd0061: exp <= 22'd4106751;
                12'd0062: exp <= 22'd4105346;
                12'd0063: exp <= 22'd4103942;
                12'd0064: exp <= 22'd4102538;
                12'd0065: exp <= 22'd4101134;
                12'd0066: exp <= 22'd4099730;
                12'd0067: exp <= 22'd4098327;
                12'd0068: exp <= 22'd4096924;
                12'd0069: exp <= 22'd4095521;
                12'd0070: exp <= 22'd4094118;
                12'd0071: exp <= 22'd4092715;
                12'd0072: exp <= 22'd4091313;
                12'd0073: exp <= 22'd4089911;
                12'd0074: exp <= 22'd4088509;
                12'd0075: exp <= 22'd4087108;
                12'd0076: exp <= 22'd4085707;
                12'd0077: exp <= 22'd4084305;
                12'd0078: exp <= 22'd4082905;
                12'd0079: exp <= 22'd4081504;
                12'd0080: exp <= 22'd4080104;
                12'd0081: exp <= 22'd4078704;
                12'd0082: exp <= 22'd4077304;
                12'd0083: exp <= 22'd4075904;
                12'd0084: exp <= 22'd4074505;
                12'd0085: exp <= 22'd4073105;
                12'd0086: exp <= 22'd4071706;
                12'd0087: exp <= 22'd4070308;
                12'd0088: exp <= 22'd4068909;
                12'd0089: exp <= 22'd4067511;
                12'd0090: exp <= 22'd4066113;
                12'd0091: exp <= 22'd4064715;
                12'd0092: exp <= 22'd4063318;
                12'd0093: exp <= 22'd4061921;
                12'd0094: exp <= 22'd4060524;
                12'd0095: exp <= 22'd4059127;
                12'd0096: exp <= 22'd4057730;
                12'd0097: exp <= 22'd4056334;
                12'd0098: exp <= 22'd4054938;
                12'd0099: exp <= 22'd4053542;
                12'd0100: exp <= 22'd4052146;
                12'd0101: exp <= 22'd4050751;
                12'd0102: exp <= 22'd4049356;
                12'd0103: exp <= 22'd4047961;
                12'd0104: exp <= 22'd4046566;
                12'd0105: exp <= 22'd4045172;
                12'd0106: exp <= 22'd4043777;
                12'd0107: exp <= 22'd4042383;
                12'd0108: exp <= 22'd4040990;
                12'd0109: exp <= 22'd4039596;
                12'd0110: exp <= 22'd4038203;
                12'd0111: exp <= 22'd4036810;
                12'd0112: exp <= 22'd4035417;
                12'd0113: exp <= 22'd4034025;
                12'd0114: exp <= 22'd4032632;
                12'd0115: exp <= 22'd4031240;
                12'd0116: exp <= 22'd4029848;
                12'd0117: exp <= 22'd4028457;
                12'd0118: exp <= 22'd4027065;
                12'd0119: exp <= 22'd4025674;
                12'd0120: exp <= 22'd4024283;
                12'd0121: exp <= 22'd4022893;
                12'd0122: exp <= 22'd4021502;
                12'd0123: exp <= 22'd4020112;
                12'd0124: exp <= 22'd4018722;
                12'd0125: exp <= 22'd4017332;
                12'd0126: exp <= 22'd4015943;
                12'd0127: exp <= 22'd4014553;
                12'd0128: exp <= 22'd4013164;
                12'd0129: exp <= 22'd4011776;
                12'd0130: exp <= 22'd4010387;
                12'd0131: exp <= 22'd4008999;
                12'd0132: exp <= 22'd4007611;
                12'd0133: exp <= 22'd4006223;
                12'd0134: exp <= 22'd4004835;
                12'd0135: exp <= 22'd4003448;
                12'd0136: exp <= 22'd4002061;
                12'd0137: exp <= 22'd4000674;
                12'd0138: exp <= 22'd3999287;
                12'd0139: exp <= 22'd3997901;
                12'd0140: exp <= 22'd3996514;
                12'd0141: exp <= 22'd3995128;
                12'd0142: exp <= 22'd3993743;
                12'd0143: exp <= 22'd3992357;
                12'd0144: exp <= 22'd3990972;
                12'd0145: exp <= 22'd3989587;
                12'd0146: exp <= 22'd3988202;
                12'd0147: exp <= 22'd3986817;
                12'd0148: exp <= 22'd3985433;
                12'd0149: exp <= 22'd3984049;
                12'd0150: exp <= 22'd3982665;
                12'd0151: exp <= 22'd3981282;
                12'd0152: exp <= 22'd3979898;
                12'd0153: exp <= 22'd3978515;
                12'd0154: exp <= 22'd3977132;
                12'd0155: exp <= 22'd3975749;
                12'd0156: exp <= 22'd3974367;
                12'd0157: exp <= 22'd3972985;
                12'd0158: exp <= 22'd3971603;
                12'd0159: exp <= 22'd3970221;
                12'd0160: exp <= 22'd3968839;
                12'd0161: exp <= 22'd3967458;
                12'd0162: exp <= 22'd3966077;
                12'd0163: exp <= 22'd3964696;
                12'd0164: exp <= 22'd3963316;
                12'd0165: exp <= 22'd3961935;
                12'd0166: exp <= 22'd3960555;
                12'd0167: exp <= 22'd3959175;
                12'd0168: exp <= 22'd3957796;
                12'd0169: exp <= 22'd3956416;
                12'd0170: exp <= 22'd3955037;
                12'd0171: exp <= 22'd3953658;
                12'd0172: exp <= 22'd3952279;
                12'd0173: exp <= 22'd3950901;
                12'd0174: exp <= 22'd3949522;
                12'd0175: exp <= 22'd3948144;
                12'd0176: exp <= 22'd3946767;
                12'd0177: exp <= 22'd3945389;
                12'd0178: exp <= 22'd3944012;
                12'd0179: exp <= 22'd3942635;
                12'd0180: exp <= 22'd3941258;
                12'd0181: exp <= 22'd3939881;
                12'd0182: exp <= 22'd3938505;
                12'd0183: exp <= 22'd3937129;
                12'd0184: exp <= 22'd3935753;
                12'd0185: exp <= 22'd3934377;
                12'd0186: exp <= 22'd3933002;
                12'd0187: exp <= 22'd3931626;
                12'd0188: exp <= 22'd3930251;
                12'd0189: exp <= 22'd3928877;
                12'd0190: exp <= 22'd3927502;
                12'd0191: exp <= 22'd3926128;
                12'd0192: exp <= 22'd3924754;
                12'd0193: exp <= 22'd3923380;
                12'd0194: exp <= 22'd3922006;
                12'd0195: exp <= 22'd3920633;
                12'd0196: exp <= 22'd3919260;
                12'd0197: exp <= 22'd3917887;
                12'd0198: exp <= 22'd3916514;
                12'd0199: exp <= 22'd3915142;
                12'd0200: exp <= 22'd3913769;
                12'd0201: exp <= 22'd3912398;
                12'd0202: exp <= 22'd3911026;
                12'd0203: exp <= 22'd3909654;
                12'd0204: exp <= 22'd3908283;
                12'd0205: exp <= 22'd3906912;
                12'd0206: exp <= 22'd3905541;
                12'd0207: exp <= 22'd3904171;
                12'd0208: exp <= 22'd3902800;
                12'd0209: exp <= 22'd3901430;
                12'd0210: exp <= 22'd3900060;
                12'd0211: exp <= 22'd3898691;
                12'd0212: exp <= 22'd3897321;
                12'd0213: exp <= 22'd3895952;
                12'd0214: exp <= 22'd3894583;
                12'd0215: exp <= 22'd3893214;
                12'd0216: exp <= 22'd3891846;
                12'd0217: exp <= 22'd3890477;
                12'd0218: exp <= 22'd3889109;
                12'd0219: exp <= 22'd3887742;
                12'd0220: exp <= 22'd3886374;
                12'd0221: exp <= 22'd3885007;
                12'd0222: exp <= 22'd3883640;
                12'd0223: exp <= 22'd3882273;
                12'd0224: exp <= 22'd3880906;
                12'd0225: exp <= 22'd3879540;
                12'd0226: exp <= 22'd3878173;
                12'd0227: exp <= 22'd3876808;
                12'd0228: exp <= 22'd3875442;
                12'd0229: exp <= 22'd3874076;
                12'd0230: exp <= 22'd3872711;
                12'd0231: exp <= 22'd3871346;
                12'd0232: exp <= 22'd3869981;
                12'd0233: exp <= 22'd3868617;
                12'd0234: exp <= 22'd3867252;
                12'd0235: exp <= 22'd3865888;
                12'd0236: exp <= 22'd3864524;
                12'd0237: exp <= 22'd3863161;
                12'd0238: exp <= 22'd3861797;
                12'd0239: exp <= 22'd3860434;
                12'd0240: exp <= 22'd3859071;
                12'd0241: exp <= 22'd3857708;
                12'd0242: exp <= 22'd3856346;
                12'd0243: exp <= 22'd3854984;
                12'd0244: exp <= 22'd3853622;
                12'd0245: exp <= 22'd3852260;
                12'd0246: exp <= 22'd3850898;
                12'd0247: exp <= 22'd3849537;
                12'd0248: exp <= 22'd3848176;
                12'd0249: exp <= 22'd3846815;
                12'd0250: exp <= 22'd3845454;
                12'd0251: exp <= 22'd3844094;
                12'd0252: exp <= 22'd3842734;
                12'd0253: exp <= 22'd3841374;
                12'd0254: exp <= 22'd3840014;
                12'd0255: exp <= 22'd3838655;
                12'd0256: exp <= 22'd3837295;
                12'd0257: exp <= 22'd3835936;
                12'd0258: exp <= 22'd3834577;
                12'd0259: exp <= 22'd3833219;
                12'd0260: exp <= 22'd3831861;
                12'd0261: exp <= 22'd3830502;
                12'd0262: exp <= 22'd3829145;
                12'd0263: exp <= 22'd3827787;
                12'd0264: exp <= 22'd3826429;
                12'd0265: exp <= 22'd3825072;
                12'd0266: exp <= 22'd3823715;
                12'd0267: exp <= 22'd3822359;
                12'd0268: exp <= 22'd3821002;
                12'd0269: exp <= 22'd3819646;
                12'd0270: exp <= 22'd3818290;
                12'd0271: exp <= 22'd3816934;
                12'd0272: exp <= 22'd3815578;
                12'd0273: exp <= 22'd3814223;
                12'd0274: exp <= 22'd3812868;
                12'd0275: exp <= 22'd3811513;
                12'd0276: exp <= 22'd3810158;
                12'd0277: exp <= 22'd3808804;
                12'd0278: exp <= 22'd3807450;
                12'd0279: exp <= 22'd3806096;
                12'd0280: exp <= 22'd3804742;
                12'd0281: exp <= 22'd3803388;
                12'd0282: exp <= 22'd3802035;
                12'd0283: exp <= 22'd3800682;
                12'd0284: exp <= 22'd3799329;
                12'd0285: exp <= 22'd3797976;
                12'd0286: exp <= 22'd3796624;
                12'd0287: exp <= 22'd3795272;
                12'd0288: exp <= 22'd3793920;
                12'd0289: exp <= 22'd3792568;
                12'd0290: exp <= 22'd3791217;
                12'd0291: exp <= 22'd3789866;
                12'd0292: exp <= 22'd3788515;
                12'd0293: exp <= 22'd3787164;
                12'd0294: exp <= 22'd3785813;
                12'd0295: exp <= 22'd3784463;
                12'd0296: exp <= 22'd3783113;
                12'd0297: exp <= 22'd3781763;
                12'd0298: exp <= 22'd3780413;
                12'd0299: exp <= 22'd3779064;
                12'd0300: exp <= 22'd3777715;
                12'd0301: exp <= 22'd3776366;
                12'd0302: exp <= 22'd3775017;
                12'd0303: exp <= 22'd3773669;
                12'd0304: exp <= 22'd3772320;
                12'd0305: exp <= 22'd3770972;
                12'd0306: exp <= 22'd3769624;
                12'd0307: exp <= 22'd3768277;
                12'd0308: exp <= 22'd3766930;
                12'd0309: exp <= 22'd3765582;
                12'd0310: exp <= 22'd3764235;
                12'd0311: exp <= 22'd3762889;
                12'd0312: exp <= 22'd3761542;
                12'd0313: exp <= 22'd3760196;
                12'd0314: exp <= 22'd3758850;
                12'd0315: exp <= 22'd3757504;
                12'd0316: exp <= 22'd3756159;
                12'd0317: exp <= 22'd3754814;
                12'd0318: exp <= 22'd3753468;
                12'd0319: exp <= 22'd3752124;
                12'd0320: exp <= 22'd3750779;
                12'd0321: exp <= 22'd3749435;
                12'd0322: exp <= 22'd3748090;
                12'd0323: exp <= 22'd3746746;
                12'd0324: exp <= 22'd3745403;
                12'd0325: exp <= 22'd3744059;
                12'd0326: exp <= 22'd3742716;
                12'd0327: exp <= 22'd3741373;
                12'd0328: exp <= 22'd3740030;
                12'd0329: exp <= 22'd3738688;
                12'd0330: exp <= 22'd3737345;
                12'd0331: exp <= 22'd3736003;
                12'd0332: exp <= 22'd3734661;
                12'd0333: exp <= 22'd3733320;
                12'd0334: exp <= 22'd3731978;
                12'd0335: exp <= 22'd3730637;
                12'd0336: exp <= 22'd3729296;
                12'd0337: exp <= 22'd3727955;
                12'd0338: exp <= 22'd3726615;
                12'd0339: exp <= 22'd3725274;
                12'd0340: exp <= 22'd3723934;
                12'd0341: exp <= 22'd3722594;
                12'd0342: exp <= 22'd3721255;
                12'd0343: exp <= 22'd3719915;
                12'd0344: exp <= 22'd3718576;
                12'd0345: exp <= 22'd3717237;
                12'd0346: exp <= 22'd3715899;
                12'd0347: exp <= 22'd3714560;
                12'd0348: exp <= 22'd3713222;
                12'd0349: exp <= 22'd3711884;
                12'd0350: exp <= 22'd3710546;
                12'd0351: exp <= 22'd3709208;
                12'd0352: exp <= 22'd3707871;
                12'd0353: exp <= 22'd3706534;
                12'd0354: exp <= 22'd3705197;
                12'd0355: exp <= 22'd3703860;
                12'd0356: exp <= 22'd3702524;
                12'd0357: exp <= 22'd3701188;
                12'd0358: exp <= 22'd3699852;
                12'd0359: exp <= 22'd3698516;
                12'd0360: exp <= 22'd3697180;
                12'd0361: exp <= 22'd3695845;
                12'd0362: exp <= 22'd3694510;
                12'd0363: exp <= 22'd3693175;
                12'd0364: exp <= 22'd3691840;
                12'd0365: exp <= 22'd3690506;
                12'd0366: exp <= 22'd3689172;
                12'd0367: exp <= 22'd3687838;
                12'd0368: exp <= 22'd3686504;
                12'd0369: exp <= 22'd3685170;
                12'd0370: exp <= 22'd3683837;
                12'd0371: exp <= 22'd3682504;
                12'd0372: exp <= 22'd3681171;
                12'd0373: exp <= 22'd3679839;
                12'd0374: exp <= 22'd3678506;
                12'd0375: exp <= 22'd3677174;
                12'd0376: exp <= 22'd3675842;
                12'd0377: exp <= 22'd3674510;
                12'd0378: exp <= 22'd3673179;
                12'd0379: exp <= 22'd3671848;
                12'd0380: exp <= 22'd3670517;
                12'd0381: exp <= 22'd3669186;
                12'd0382: exp <= 22'd3667855;
                12'd0383: exp <= 22'd3666525;
                12'd0384: exp <= 22'd3665195;
                12'd0385: exp <= 22'd3663865;
                12'd0386: exp <= 22'd3662535;
                12'd0387: exp <= 22'd3661206;
                12'd0388: exp <= 22'd3659876;
                12'd0389: exp <= 22'd3658547;
                12'd0390: exp <= 22'd3657219;
                12'd0391: exp <= 22'd3655890;
                12'd0392: exp <= 22'd3654562;
                12'd0393: exp <= 22'd3653234;
                12'd0394: exp <= 22'd3651906;
                12'd0395: exp <= 22'd3650578;
                12'd0396: exp <= 22'd3649251;
                12'd0397: exp <= 22'd3647923;
                12'd0398: exp <= 22'd3646596;
                12'd0399: exp <= 22'd3645270;
                12'd0400: exp <= 22'd3643943;
                12'd0401: exp <= 22'd3642617;
                12'd0402: exp <= 22'd3641291;
                12'd0403: exp <= 22'd3639965;
                12'd0404: exp <= 22'd3638639;
                12'd0405: exp <= 22'd3637314;
                12'd0406: exp <= 22'd3635988;
                12'd0407: exp <= 22'd3634664;
                12'd0408: exp <= 22'd3633339;
                12'd0409: exp <= 22'd3632014;
                12'd0410: exp <= 22'd3630690;
                12'd0411: exp <= 22'd3629366;
                12'd0412: exp <= 22'd3628042;
                12'd0413: exp <= 22'd3626718;
                12'd0414: exp <= 22'd3625395;
                12'd0415: exp <= 22'd3624072;
                12'd0416: exp <= 22'd3622749;
                12'd0417: exp <= 22'd3621426;
                12'd0418: exp <= 22'd3620104;
                12'd0419: exp <= 22'd3618781;
                12'd0420: exp <= 22'd3617459;
                12'd0421: exp <= 22'd3616137;
                12'd0422: exp <= 22'd3614816;
                12'd0423: exp <= 22'd3613494;
                12'd0424: exp <= 22'd3612173;
                12'd0425: exp <= 22'd3610852;
                12'd0426: exp <= 22'd3609532;
                12'd0427: exp <= 22'd3608211;
                12'd0428: exp <= 22'd3606891;
                12'd0429: exp <= 22'd3605571;
                12'd0430: exp <= 22'd3604251;
                12'd0431: exp <= 22'd3602931;
                12'd0432: exp <= 22'd3601612;
                12'd0433: exp <= 22'd3600293;
                12'd0434: exp <= 22'd3598974;
                12'd0435: exp <= 22'd3597655;
                12'd0436: exp <= 22'd3596337;
                12'd0437: exp <= 22'd3595018;
                12'd0438: exp <= 22'd3593700;
                12'd0439: exp <= 22'd3592383;
                12'd0440: exp <= 22'd3591065;
                12'd0441: exp <= 22'd3589748;
                12'd0442: exp <= 22'd3588430;
                12'd0443: exp <= 22'd3587114;
                12'd0444: exp <= 22'd3585797;
                12'd0445: exp <= 22'd3584480;
                12'd0446: exp <= 22'd3583164;
                12'd0447: exp <= 22'd3581848;
                12'd0448: exp <= 22'd3580532;
                12'd0449: exp <= 22'd3579217;
                12'd0450: exp <= 22'd3577901;
                12'd0451: exp <= 22'd3576586;
                12'd0452: exp <= 22'd3575271;
                12'd0453: exp <= 22'd3573957;
                12'd0454: exp <= 22'd3572642;
                12'd0455: exp <= 22'd3571328;
                12'd0456: exp <= 22'd3570014;
                12'd0457: exp <= 22'd3568700;
                12'd0458: exp <= 22'd3567386;
                12'd0459: exp <= 22'd3566073;
                12'd0460: exp <= 22'd3564760;
                12'd0461: exp <= 22'd3563447;
                12'd0462: exp <= 22'd3562134;
                12'd0463: exp <= 22'd3560822;
                12'd0464: exp <= 22'd3559510;
                12'd0465: exp <= 22'd3558197;
                12'd0466: exp <= 22'd3556886;
                12'd0467: exp <= 22'd3555574;
                12'd0468: exp <= 22'd3554263;
                12'd0469: exp <= 22'd3552952;
                12'd0470: exp <= 22'd3551641;
                12'd0471: exp <= 22'd3550330;
                12'd0472: exp <= 22'd3549019;
                12'd0473: exp <= 22'd3547709;
                12'd0474: exp <= 22'd3546399;
                12'd0475: exp <= 22'd3545089;
                12'd0476: exp <= 22'd3543780;
                12'd0477: exp <= 22'd3542470;
                12'd0478: exp <= 22'd3541161;
                12'd0479: exp <= 22'd3539852;
                12'd0480: exp <= 22'd3538544;
                12'd0481: exp <= 22'd3537235;
                12'd0482: exp <= 22'd3535927;
                12'd0483: exp <= 22'd3534619;
                12'd0484: exp <= 22'd3533311;
                12'd0485: exp <= 22'd3532003;
                12'd0486: exp <= 22'd3530696;
                12'd0487: exp <= 22'd3529389;
                12'd0488: exp <= 22'd3528082;
                12'd0489: exp <= 22'd3526775;
                12'd0490: exp <= 22'd3525469;
                12'd0491: exp <= 22'd3524163;
                12'd0492: exp <= 22'd3522856;
                12'd0493: exp <= 22'd3521551;
                12'd0494: exp <= 22'd3520245;
                12'd0495: exp <= 22'd3518940;
                12'd0496: exp <= 22'd3517634;
                12'd0497: exp <= 22'd3516330;
                12'd0498: exp <= 22'd3515025;
                12'd0499: exp <= 22'd3513720;
                12'd0500: exp <= 22'd3512416;
                12'd0501: exp <= 22'd3511112;
                12'd0502: exp <= 22'd3509808;
                12'd0503: exp <= 22'd3508504;
                12'd0504: exp <= 22'd3507201;
                12'd0505: exp <= 22'd3505898;
                12'd0506: exp <= 22'd3504595;
                12'd0507: exp <= 22'd3503292;
                12'd0508: exp <= 22'd3501990;
                12'd0509: exp <= 22'd3500687;
                12'd0510: exp <= 22'd3499385;
                12'd0511: exp <= 22'd3498083;
                12'd0512: exp <= 22'd3496782;
                12'd0513: exp <= 22'd3495480;
                12'd0514: exp <= 22'd3494179;
                12'd0515: exp <= 22'd3492878;
                12'd0516: exp <= 22'd3491577;
                12'd0517: exp <= 22'd3490277;
                12'd0518: exp <= 22'd3488977;
                12'd0519: exp <= 22'd3487677;
                12'd0520: exp <= 22'd3486377;
                12'd0521: exp <= 22'd3485077;
                12'd0522: exp <= 22'd3483778;
                12'd0523: exp <= 22'd3482478;
                12'd0524: exp <= 22'd3481179;
                12'd0525: exp <= 22'd3479881;
                12'd0526: exp <= 22'd3478582;
                12'd0527: exp <= 22'd3477284;
                12'd0528: exp <= 22'd3475986;
                12'd0529: exp <= 22'd3474688;
                12'd0530: exp <= 22'd3473390;
                12'd0531: exp <= 22'd3472093;
                12'd0532: exp <= 22'd3470795;
                12'd0533: exp <= 22'd3469498;
                12'd0534: exp <= 22'd3468201;
                12'd0535: exp <= 22'd3466905;
                12'd0536: exp <= 22'd3465609;
                12'd0537: exp <= 22'd3464312;
                12'd0538: exp <= 22'd3463016;
                12'd0539: exp <= 22'd3461721;
                12'd0540: exp <= 22'd3460425;
                12'd0541: exp <= 22'd3459130;
                12'd0542: exp <= 22'd3457835;
                12'd0543: exp <= 22'd3456540;
                12'd0544: exp <= 22'd3455246;
                12'd0545: exp <= 22'd3453951;
                12'd0546: exp <= 22'd3452657;
                12'd0547: exp <= 22'd3451363;
                12'd0548: exp <= 22'd3450069;
                12'd0549: exp <= 22'd3448776;
                12'd0550: exp <= 22'd3447482;
                12'd0551: exp <= 22'd3446189;
                12'd0552: exp <= 22'd3444897;
                12'd0553: exp <= 22'd3443604;
                12'd0554: exp <= 22'd3442311;
                12'd0555: exp <= 22'd3441019;
                12'd0556: exp <= 22'd3439727;
                12'd0557: exp <= 22'd3438436;
                12'd0558: exp <= 22'd3437144;
                12'd0559: exp <= 22'd3435853;
                12'd0560: exp <= 22'd3434562;
                12'd0561: exp <= 22'd3433271;
                12'd0562: exp <= 22'd3431980;
                12'd0563: exp <= 22'd3430690;
                12'd0564: exp <= 22'd3429399;
                12'd0565: exp <= 22'd3428109;
                12'd0566: exp <= 22'd3426820;
                12'd0567: exp <= 22'd3425530;
                12'd0568: exp <= 22'd3424241;
                12'd0569: exp <= 22'd3422951;
                12'd0570: exp <= 22'd3421663;
                12'd0571: exp <= 22'd3420374;
                12'd0572: exp <= 22'd3419085;
                12'd0573: exp <= 22'd3417797;
                12'd0574: exp <= 22'd3416509;
                12'd0575: exp <= 22'd3415221;
                12'd0576: exp <= 22'd3413934;
                12'd0577: exp <= 22'd3412646;
                12'd0578: exp <= 22'd3411359;
                12'd0579: exp <= 22'd3410072;
                12'd0580: exp <= 22'd3408785;
                12'd0581: exp <= 22'd3407499;
                12'd0582: exp <= 22'd3406212;
                12'd0583: exp <= 22'd3404926;
                12'd0584: exp <= 22'd3403640;
                12'd0585: exp <= 22'd3402355;
                12'd0586: exp <= 22'd3401069;
                12'd0587: exp <= 22'd3399784;
                12'd0588: exp <= 22'd3398499;
                12'd0589: exp <= 22'd3397214;
                12'd0590: exp <= 22'd3395930;
                12'd0591: exp <= 22'd3394645;
                12'd0592: exp <= 22'd3393361;
                12'd0593: exp <= 22'd3392077;
                12'd0594: exp <= 22'd3390794;
                12'd0595: exp <= 22'd3389510;
                12'd0596: exp <= 22'd3388227;
                12'd0597: exp <= 22'd3386944;
                12'd0598: exp <= 22'd3385661;
                12'd0599: exp <= 22'd3384378;
                12'd0600: exp <= 22'd3383096;
                12'd0601: exp <= 22'd3381814;
                12'd0602: exp <= 22'd3380532;
                12'd0603: exp <= 22'd3379250;
                12'd0604: exp <= 22'd3377969;
                12'd0605: exp <= 22'd3376687;
                12'd0606: exp <= 22'd3375406;
                12'd0607: exp <= 22'd3374125;
                12'd0608: exp <= 22'd3372845;
                12'd0609: exp <= 22'd3371564;
                12'd0610: exp <= 22'd3370284;
                12'd0611: exp <= 22'd3369004;
                12'd0612: exp <= 22'd3367724;
                12'd0613: exp <= 22'd3366445;
                12'd0614: exp <= 22'd3365165;
                12'd0615: exp <= 22'd3363886;
                12'd0616: exp <= 22'd3362607;
                12'd0617: exp <= 22'd3361328;
                12'd0618: exp <= 22'd3360050;
                12'd0619: exp <= 22'd3358772;
                12'd0620: exp <= 22'd3357494;
                12'd0621: exp <= 22'd3356216;
                12'd0622: exp <= 22'd3354938;
                12'd0623: exp <= 22'd3353661;
                12'd0624: exp <= 22'd3352384;
                12'd0625: exp <= 22'd3351107;
                12'd0626: exp <= 22'd3349830;
                12'd0627: exp <= 22'd3348553;
                12'd0628: exp <= 22'd3347277;
                12'd0629: exp <= 22'd3346001;
                12'd0630: exp <= 22'd3344725;
                12'd0631: exp <= 22'd3343449;
                12'd0632: exp <= 22'd3342174;
                12'd0633: exp <= 22'd3340898;
                12'd0634: exp <= 22'd3339623;
                12'd0635: exp <= 22'd3338349;
                12'd0636: exp <= 22'd3337074;
                12'd0637: exp <= 22'd3335800;
                12'd0638: exp <= 22'd3334525;
                12'd0639: exp <= 22'd3333251;
                12'd0640: exp <= 22'd3331978;
                12'd0641: exp <= 22'd3330704;
                12'd0642: exp <= 22'd3329431;
                12'd0643: exp <= 22'd3328158;
                12'd0644: exp <= 22'd3326885;
                12'd0645: exp <= 22'd3325612;
                12'd0646: exp <= 22'd3324340;
                12'd0647: exp <= 22'd3323068;
                12'd0648: exp <= 22'd3321795;
                12'd0649: exp <= 22'd3320524;
                12'd0650: exp <= 22'd3319252;
                12'd0651: exp <= 22'd3317981;
                12'd0652: exp <= 22'd3316710;
                12'd0653: exp <= 22'd3315439;
                12'd0654: exp <= 22'd3314168;
                12'd0655: exp <= 22'd3312897;
                12'd0656: exp <= 22'd3311627;
                12'd0657: exp <= 22'd3310357;
                12'd0658: exp <= 22'd3309087;
                12'd0659: exp <= 22'd3307817;
                12'd0660: exp <= 22'd3306548;
                12'd0661: exp <= 22'd3305279;
                12'd0662: exp <= 22'd3304010;
                12'd0663: exp <= 22'd3302741;
                12'd0664: exp <= 22'd3301472;
                12'd0665: exp <= 22'd3300204;
                12'd0666: exp <= 22'd3298936;
                12'd0667: exp <= 22'd3297668;
                12'd0668: exp <= 22'd3296400;
                12'd0669: exp <= 22'd3295133;
                12'd0670: exp <= 22'd3293865;
                12'd0671: exp <= 22'd3292598;
                12'd0672: exp <= 22'd3291331;
                12'd0673: exp <= 22'd3290065;
                12'd0674: exp <= 22'd3288798;
                12'd0675: exp <= 22'd3287532;
                12'd0676: exp <= 22'd3286266;
                12'd0677: exp <= 22'd3285000;
                12'd0678: exp <= 22'd3283735;
                12'd0679: exp <= 22'd3282469;
                12'd0680: exp <= 22'd3281204;
                12'd0681: exp <= 22'd3279939;
                12'd0682: exp <= 22'd3278675;
                12'd0683: exp <= 22'd3277410;
                12'd0684: exp <= 22'd3276146;
                12'd0685: exp <= 22'd3274882;
                12'd0686: exp <= 22'd3273618;
                12'd0687: exp <= 22'd3272354;
                12'd0688: exp <= 22'd3271091;
                12'd0689: exp <= 22'd3269827;
                12'd0690: exp <= 22'd3268564;
                12'd0691: exp <= 22'd3267302;
                12'd0692: exp <= 22'd3266039;
                12'd0693: exp <= 22'd3264777;
                12'd0694: exp <= 22'd3263515;
                12'd0695: exp <= 22'd3262253;
                12'd0696: exp <= 22'd3260991;
                12'd0697: exp <= 22'd3259729;
                12'd0698: exp <= 22'd3258468;
                12'd0699: exp <= 22'd3257207;
                12'd0700: exp <= 22'd3255946;
                12'd0701: exp <= 22'd3254685;
                12'd0702: exp <= 22'd3253425;
                12'd0703: exp <= 22'd3252165;
                12'd0704: exp <= 22'd3250905;
                12'd0705: exp <= 22'd3249645;
                12'd0706: exp <= 22'd3248385;
                12'd0707: exp <= 22'd3247126;
                12'd0708: exp <= 22'd3245867;
                12'd0709: exp <= 22'd3244608;
                12'd0710: exp <= 22'd3243349;
                12'd0711: exp <= 22'd3242090;
                12'd0712: exp <= 22'd3240832;
                12'd0713: exp <= 22'd3239574;
                12'd0714: exp <= 22'd3238316;
                12'd0715: exp <= 22'd3237058;
                12'd0716: exp <= 22'd3235801;
                12'd0717: exp <= 22'd3234544;
                12'd0718: exp <= 22'd3233287;
                12'd0719: exp <= 22'd3232030;
                12'd0720: exp <= 22'd3230773;
                12'd0721: exp <= 22'd3229517;
                12'd0722: exp <= 22'd3228261;
                12'd0723: exp <= 22'd3227005;
                12'd0724: exp <= 22'd3225749;
                12'd0725: exp <= 22'd3224493;
                12'd0726: exp <= 22'd3223238;
                12'd0727: exp <= 22'd3221983;
                12'd0728: exp <= 22'd3220728;
                12'd0729: exp <= 22'd3219473;
                12'd0730: exp <= 22'd3218219;
                12'd0731: exp <= 22'd3216965;
                12'd0732: exp <= 22'd3215710;
                12'd0733: exp <= 22'd3214457;
                12'd0734: exp <= 22'd3213203;
                12'd0735: exp <= 22'd3211949;
                12'd0736: exp <= 22'd3210696;
                12'd0737: exp <= 22'd3209443;
                12'd0738: exp <= 22'd3208190;
                12'd0739: exp <= 22'd3206938;
                12'd0740: exp <= 22'd3205686;
                12'd0741: exp <= 22'd3204433;
                12'd0742: exp <= 22'd3203181;
                12'd0743: exp <= 22'd3201930;
                12'd0744: exp <= 22'd3200678;
                12'd0745: exp <= 22'd3199427;
                12'd0746: exp <= 22'd3198176;
                12'd0747: exp <= 22'd3196925;
                12'd0748: exp <= 22'd3195674;
                12'd0749: exp <= 22'd3194424;
                12'd0750: exp <= 22'd3193173;
                12'd0751: exp <= 22'd3191923;
                12'd0752: exp <= 22'd3190674;
                12'd0753: exp <= 22'd3189424;
                12'd0754: exp <= 22'd3188175;
                12'd0755: exp <= 22'd3186925;
                12'd0756: exp <= 22'd3185676;
                12'd0757: exp <= 22'd3184428;
                12'd0758: exp <= 22'd3183179;
                12'd0759: exp <= 22'd3181931;
                12'd0760: exp <= 22'd3180683;
                12'd0761: exp <= 22'd3179435;
                12'd0762: exp <= 22'd3178187;
                12'd0763: exp <= 22'd3176939;
                12'd0764: exp <= 22'd3175692;
                12'd0765: exp <= 22'd3174445;
                12'd0766: exp <= 22'd3173198;
                12'd0767: exp <= 22'd3171951;
                12'd0768: exp <= 22'd3170705;
                12'd0769: exp <= 22'd3169459;
                12'd0770: exp <= 22'd3168213;
                12'd0771: exp <= 22'd3166967;
                12'd0772: exp <= 22'd3165721;
                12'd0773: exp <= 22'd3164476;
                12'd0774: exp <= 22'd3163231;
                12'd0775: exp <= 22'd3161986;
                12'd0776: exp <= 22'd3160741;
                12'd0777: exp <= 22'd3159496;
                12'd0778: exp <= 22'd3158252;
                12'd0779: exp <= 22'd3157008;
                12'd0780: exp <= 22'd3155764;
                12'd0781: exp <= 22'd3154520;
                12'd0782: exp <= 22'd3153277;
                12'd0783: exp <= 22'd3152034;
                12'd0784: exp <= 22'd3150790;
                12'd0785: exp <= 22'd3149548;
                12'd0786: exp <= 22'd3148305;
                12'd0787: exp <= 22'd3147062;
                12'd0788: exp <= 22'd3145820;
                12'd0789: exp <= 22'd3144578;
                12'd0790: exp <= 22'd3143336;
                12'd0791: exp <= 22'd3142095;
                12'd0792: exp <= 22'd3140853;
                12'd0793: exp <= 22'd3139612;
                12'd0794: exp <= 22'd3138371;
                12'd0795: exp <= 22'd3137130;
                12'd0796: exp <= 22'd3135890;
                12'd0797: exp <= 22'd3134650;
                12'd0798: exp <= 22'd3133409;
                12'd0799: exp <= 22'd3132169;
                12'd0800: exp <= 22'd3130930;
                12'd0801: exp <= 22'd3129690;
                12'd0802: exp <= 22'd3128451;
                12'd0803: exp <= 22'd3127212;
                12'd0804: exp <= 22'd3125973;
                12'd0805: exp <= 22'd3124734;
                12'd0806: exp <= 22'd3123496;
                12'd0807: exp <= 22'd3122258;
                12'd0808: exp <= 22'd3121020;
                12'd0809: exp <= 22'd3119782;
                12'd0810: exp <= 22'd3118544;
                12'd0811: exp <= 22'd3117307;
                12'd0812: exp <= 22'd3116069;
                12'd0813: exp <= 22'd3114832;
                12'd0814: exp <= 22'd3113596;
                12'd0815: exp <= 22'd3112359;
                12'd0816: exp <= 22'd3111123;
                12'd0817: exp <= 22'd3109887;
                12'd0818: exp <= 22'd3108651;
                12'd0819: exp <= 22'd3107415;
                12'd0820: exp <= 22'd3106179;
                12'd0821: exp <= 22'd3104944;
                12'd0822: exp <= 22'd3103709;
                12'd0823: exp <= 22'd3102474;
                12'd0824: exp <= 22'd3101239;
                12'd0825: exp <= 22'd3100005;
                12'd0826: exp <= 22'd3098771;
                12'd0827: exp <= 22'd3097536;
                12'd0828: exp <= 22'd3096303;
                12'd0829: exp <= 22'd3095069;
                12'd0830: exp <= 22'd3093835;
                12'd0831: exp <= 22'd3092602;
                12'd0832: exp <= 22'd3091369;
                12'd0833: exp <= 22'd3090136;
                12'd0834: exp <= 22'd3088904;
                12'd0835: exp <= 22'd3087671;
                12'd0836: exp <= 22'd3086439;
                12'd0837: exp <= 22'd3085207;
                12'd0838: exp <= 22'd3083975;
                12'd0839: exp <= 22'd3082744;
                12'd0840: exp <= 22'd3081513;
                12'd0841: exp <= 22'd3080281;
                12'd0842: exp <= 22'd3079050;
                12'd0843: exp <= 22'd3077820;
                12'd0844: exp <= 22'd3076589;
                12'd0845: exp <= 22'd3075359;
                12'd0846: exp <= 22'd3074129;
                12'd0847: exp <= 22'd3072899;
                12'd0848: exp <= 22'd3071669;
                12'd0849: exp <= 22'd3070440;
                12'd0850: exp <= 22'd3069210;
                12'd0851: exp <= 22'd3067981;
                12'd0852: exp <= 22'd3066752;
                12'd0853: exp <= 22'd3065524;
                12'd0854: exp <= 22'd3064295;
                12'd0855: exp <= 22'd3063067;
                12'd0856: exp <= 22'd3061839;
                12'd0857: exp <= 22'd3060611;
                12'd0858: exp <= 22'd3059384;
                12'd0859: exp <= 22'd3058156;
                12'd0860: exp <= 22'd3056929;
                12'd0861: exp <= 22'd3055702;
                12'd0862: exp <= 22'd3054475;
                12'd0863: exp <= 22'd3053249;
                12'd0864: exp <= 22'd3052022;
                12'd0865: exp <= 22'd3050796;
                12'd0866: exp <= 22'd3049570;
                12'd0867: exp <= 22'd3048345;
                12'd0868: exp <= 22'd3047119;
                12'd0869: exp <= 22'd3045894;
                12'd0870: exp <= 22'd3044669;
                12'd0871: exp <= 22'd3043444;
                12'd0872: exp <= 22'd3042219;
                12'd0873: exp <= 22'd3040994;
                12'd0874: exp <= 22'd3039770;
                12'd0875: exp <= 22'd3038546;
                12'd0876: exp <= 22'd3037322;
                12'd0877: exp <= 22'd3036099;
                12'd0878: exp <= 22'd3034875;
                12'd0879: exp <= 22'd3033652;
                12'd0880: exp <= 22'd3032429;
                12'd0881: exp <= 22'd3031206;
                12'd0882: exp <= 22'd3029983;
                12'd0883: exp <= 22'd3028761;
                12'd0884: exp <= 22'd3027539;
                12'd0885: exp <= 22'd3026317;
                12'd0886: exp <= 22'd3025095;
                12'd0887: exp <= 22'd3023873;
                12'd0888: exp <= 22'd3022652;
                12'd0889: exp <= 22'd3021431;
                12'd0890: exp <= 22'd3020210;
                12'd0891: exp <= 22'd3018989;
                12'd0892: exp <= 22'd3017768;
                12'd0893: exp <= 22'd3016548;
                12'd0894: exp <= 22'd3015328;
                12'd0895: exp <= 22'd3014108;
                12'd0896: exp <= 22'd3012888;
                12'd0897: exp <= 22'd3011669;
                12'd0898: exp <= 22'd3010449;
                12'd0899: exp <= 22'd3009230;
                12'd0900: exp <= 22'd3008011;
                12'd0901: exp <= 22'd3006792;
                12'd0902: exp <= 22'd3005574;
                12'd0903: exp <= 22'd3004356;
                12'd0904: exp <= 22'd3003138;
                12'd0905: exp <= 22'd3001920;
                12'd0906: exp <= 22'd3000702;
                12'd0907: exp <= 22'd2999484;
                12'd0908: exp <= 22'd2998267;
                12'd0909: exp <= 22'd2997050;
                12'd0910: exp <= 22'd2995833;
                12'd0911: exp <= 22'd2994617;
                12'd0912: exp <= 22'd2993400;
                12'd0913: exp <= 22'd2992184;
                12'd0914: exp <= 22'd2990968;
                12'd0915: exp <= 22'd2989752;
                12'd0916: exp <= 22'd2988536;
                12'd0917: exp <= 22'd2987321;
                12'd0918: exp <= 22'd2986106;
                12'd0919: exp <= 22'd2984891;
                12'd0920: exp <= 22'd2983676;
                12'd0921: exp <= 22'd2982461;
                12'd0922: exp <= 22'd2981247;
                12'd0923: exp <= 22'd2980033;
                12'd0924: exp <= 22'd2978819;
                12'd0925: exp <= 22'd2977605;
                12'd0926: exp <= 22'd2976392;
                12'd0927: exp <= 22'd2975178;
                12'd0928: exp <= 22'd2973965;
                12'd0929: exp <= 22'd2972752;
                12'd0930: exp <= 22'd2971539;
                12'd0931: exp <= 22'd2970327;
                12'd0932: exp <= 22'd2969114;
                12'd0933: exp <= 22'd2967902;
                12'd0934: exp <= 22'd2966690;
                12'd0935: exp <= 22'd2965479;
                12'd0936: exp <= 22'd2964267;
                12'd0937: exp <= 22'd2963056;
                12'd0938: exp <= 22'd2961845;
                12'd0939: exp <= 22'd2960634;
                12'd0940: exp <= 22'd2959423;
                12'd0941: exp <= 22'd2958213;
                12'd0942: exp <= 22'd2957002;
                12'd0943: exp <= 22'd2955792;
                12'd0944: exp <= 22'd2954582;
                12'd0945: exp <= 22'd2953373;
                12'd0946: exp <= 22'd2952163;
                12'd0947: exp <= 22'd2950954;
                12'd0948: exp <= 22'd2949745;
                12'd0949: exp <= 22'd2948536;
                12'd0950: exp <= 22'd2947328;
                12'd0951: exp <= 22'd2946119;
                12'd0952: exp <= 22'd2944911;
                12'd0953: exp <= 22'd2943703;
                12'd0954: exp <= 22'd2942495;
                12'd0955: exp <= 22'd2941287;
                12'd0956: exp <= 22'd2940080;
                12'd0957: exp <= 22'd2938873;
                12'd0958: exp <= 22'd2937666;
                12'd0959: exp <= 22'd2936459;
                12'd0960: exp <= 22'd2935252;
                12'd0961: exp <= 22'd2934046;
                12'd0962: exp <= 22'd2932840;
                12'd0963: exp <= 22'd2931634;
                12'd0964: exp <= 22'd2930428;
                12'd0965: exp <= 22'd2929222;
                12'd0966: exp <= 22'd2928017;
                12'd0967: exp <= 22'd2926812;
                12'd0968: exp <= 22'd2925607;
                12'd0969: exp <= 22'd2924402;
                12'd0970: exp <= 22'd2923197;
                12'd0971: exp <= 22'd2921993;
                12'd0972: exp <= 22'd2920789;
                12'd0973: exp <= 22'd2919585;
                12'd0974: exp <= 22'd2918381;
                12'd0975: exp <= 22'd2917178;
                12'd0976: exp <= 22'd2915974;
                12'd0977: exp <= 22'd2914771;
                12'd0978: exp <= 22'd2913568;
                12'd0979: exp <= 22'd2912366;
                12'd0980: exp <= 22'd2911163;
                12'd0981: exp <= 22'd2909961;
                12'd0982: exp <= 22'd2908759;
                12'd0983: exp <= 22'd2907557;
                12'd0984: exp <= 22'd2906355;
                12'd0985: exp <= 22'd2905153;
                12'd0986: exp <= 22'd2903952;
                12'd0987: exp <= 22'd2902751;
                12'd0988: exp <= 22'd2901550;
                12'd0989: exp <= 22'd2900349;
                12'd0990: exp <= 22'd2899149;
                12'd0991: exp <= 22'd2897949;
                12'd0992: exp <= 22'd2896749;
                12'd0993: exp <= 22'd2895549;
                12'd0994: exp <= 22'd2894349;
                12'd0995: exp <= 22'd2893150;
                12'd0996: exp <= 22'd2891950;
                12'd0997: exp <= 22'd2890751;
                12'd0998: exp <= 22'd2889552;
                12'd0999: exp <= 22'd2888354;
                12'd1000: exp <= 22'd2887155;
                12'd1001: exp <= 22'd2885957;
                12'd1002: exp <= 22'd2884759;
                12'd1003: exp <= 22'd2883561;
                12'd1004: exp <= 22'd2882363;
                12'd1005: exp <= 22'd2881166;
                12'd1006: exp <= 22'd2879969;
                12'd1007: exp <= 22'd2878772;
                12'd1008: exp <= 22'd2877575;
                12'd1009: exp <= 22'd2876378;
                12'd1010: exp <= 22'd2875182;
                12'd1011: exp <= 22'd2873985;
                12'd1012: exp <= 22'd2872789;
                12'd1013: exp <= 22'd2871594;
                12'd1014: exp <= 22'd2870398;
                12'd1015: exp <= 22'd2869203;
                12'd1016: exp <= 22'd2868007;
                12'd1017: exp <= 22'd2866812;
                12'd1018: exp <= 22'd2865617;
                12'd1019: exp <= 22'd2864423;
                12'd1020: exp <= 22'd2863228;
                12'd1021: exp <= 22'd2862034;
                12'd1022: exp <= 22'd2860840;
                12'd1023: exp <= 22'd2859646;
                12'd1024: exp <= 22'd2858453;
                12'd1025: exp <= 22'd2857259;
                12'd1026: exp <= 22'd2856066;
                12'd1027: exp <= 22'd2854873;
                12'd1028: exp <= 22'd2853680;
                12'd1029: exp <= 22'd2852488;
                12'd1030: exp <= 22'd2851295;
                12'd1031: exp <= 22'd2850103;
                12'd1032: exp <= 22'd2848911;
                12'd1033: exp <= 22'd2847719;
                12'd1034: exp <= 22'd2846528;
                12'd1035: exp <= 22'd2845336;
                12'd1036: exp <= 22'd2844145;
                12'd1037: exp <= 22'd2842954;
                12'd1038: exp <= 22'd2841763;
                12'd1039: exp <= 22'd2840573;
                12'd1040: exp <= 22'd2839383;
                12'd1041: exp <= 22'd2838192;
                12'd1042: exp <= 22'd2837002;
                12'd1043: exp <= 22'd2835813;
                12'd1044: exp <= 22'd2834623;
                12'd1045: exp <= 22'd2833434;
                12'd1046: exp <= 22'd2832244;
                12'd1047: exp <= 22'd2831056;
                12'd1048: exp <= 22'd2829867;
                12'd1049: exp <= 22'd2828678;
                12'd1050: exp <= 22'd2827490;
                12'd1051: exp <= 22'd2826302;
                12'd1052: exp <= 22'd2825114;
                12'd1053: exp <= 22'd2823926;
                12'd1054: exp <= 22'd2822738;
                12'd1055: exp <= 22'd2821551;
                12'd1056: exp <= 22'd2820364;
                12'd1057: exp <= 22'd2819177;
                12'd1058: exp <= 22'd2817990;
                12'd1059: exp <= 22'd2816804;
                12'd1060: exp <= 22'd2815617;
                12'd1061: exp <= 22'd2814431;
                12'd1062: exp <= 22'd2813245;
                12'd1063: exp <= 22'd2812059;
                12'd1064: exp <= 22'd2810874;
                12'd1065: exp <= 22'd2809688;
                12'd1066: exp <= 22'd2808503;
                12'd1067: exp <= 22'd2807318;
                12'd1068: exp <= 22'd2806134;
                12'd1069: exp <= 22'd2804949;
                12'd1070: exp <= 22'd2803765;
                12'd1071: exp <= 22'd2802581;
                12'd1072: exp <= 22'd2801397;
                12'd1073: exp <= 22'd2800213;
                12'd1074: exp <= 22'd2799029;
                12'd1075: exp <= 22'd2797846;
                12'd1076: exp <= 22'd2796663;
                12'd1077: exp <= 22'd2795480;
                12'd1078: exp <= 22'd2794297;
                12'd1079: exp <= 22'd2793115;
                12'd1080: exp <= 22'd2791932;
                12'd1081: exp <= 22'd2790750;
                12'd1082: exp <= 22'd2789568;
                12'd1083: exp <= 22'd2788386;
                12'd1084: exp <= 22'd2787205;
                12'd1085: exp <= 22'd2786023;
                12'd1086: exp <= 22'd2784842;
                12'd1087: exp <= 22'd2783661;
                12'd1088: exp <= 22'd2782481;
                12'd1089: exp <= 22'd2781300;
                12'd1090: exp <= 22'd2780120;
                12'd1091: exp <= 22'd2778940;
                12'd1092: exp <= 22'd2777760;
                12'd1093: exp <= 22'd2776580;
                12'd1094: exp <= 22'd2775400;
                12'd1095: exp <= 22'd2774221;
                12'd1096: exp <= 22'd2773042;
                12'd1097: exp <= 22'd2771863;
                12'd1098: exp <= 22'd2770684;
                12'd1099: exp <= 22'd2769506;
                12'd1100: exp <= 22'd2768327;
                12'd1101: exp <= 22'd2767149;
                12'd1102: exp <= 22'd2765971;
                12'd1103: exp <= 22'd2764793;
                12'd1104: exp <= 22'd2763616;
                12'd1105: exp <= 22'd2762438;
                12'd1106: exp <= 22'd2761261;
                12'd1107: exp <= 22'd2760084;
                12'd1108: exp <= 22'd2758908;
                12'd1109: exp <= 22'd2757731;
                12'd1110: exp <= 22'd2756555;
                12'd1111: exp <= 22'd2755378;
                12'd1112: exp <= 22'd2754202;
                12'd1113: exp <= 22'd2753027;
                12'd1114: exp <= 22'd2751851;
                12'd1115: exp <= 22'd2750676;
                12'd1116: exp <= 22'd2749501;
                12'd1117: exp <= 22'd2748326;
                12'd1118: exp <= 22'd2747151;
                12'd1119: exp <= 22'd2745976;
                12'd1120: exp <= 22'd2744802;
                12'd1121: exp <= 22'd2743628;
                12'd1122: exp <= 22'd2742454;
                12'd1123: exp <= 22'd2741280;
                12'd1124: exp <= 22'd2740106;
                12'd1125: exp <= 22'd2738933;
                12'd1126: exp <= 22'd2737760;
                12'd1127: exp <= 22'd2736587;
                12'd1128: exp <= 22'd2735414;
                12'd1129: exp <= 22'd2734242;
                12'd1130: exp <= 22'd2733069;
                12'd1131: exp <= 22'd2731897;
                12'd1132: exp <= 22'd2730725;
                12'd1133: exp <= 22'd2729553;
                12'd1134: exp <= 22'd2728382;
                12'd1135: exp <= 22'd2727210;
                12'd1136: exp <= 22'd2726039;
                12'd1137: exp <= 22'd2724868;
                12'd1138: exp <= 22'd2723697;
                12'd1139: exp <= 22'd2722527;
                12'd1140: exp <= 22'd2721356;
                12'd1141: exp <= 22'd2720186;
                12'd1142: exp <= 22'd2719016;
                12'd1143: exp <= 22'd2717846;
                12'd1144: exp <= 22'd2716677;
                12'd1145: exp <= 22'd2715507;
                12'd1146: exp <= 22'd2714338;
                12'd1147: exp <= 22'd2713169;
                12'd1148: exp <= 22'd2712000;
                12'd1149: exp <= 22'd2710831;
                12'd1150: exp <= 22'd2709663;
                12'd1151: exp <= 22'd2708495;
                12'd1152: exp <= 22'd2707327;
                12'd1153: exp <= 22'd2706159;
                12'd1154: exp <= 22'd2704991;
                12'd1155: exp <= 22'd2703824;
                12'd1156: exp <= 22'd2702657;
                12'd1157: exp <= 22'd2701490;
                12'd1158: exp <= 22'd2700323;
                12'd1159: exp <= 22'd2699156;
                12'd1160: exp <= 22'd2697990;
                12'd1161: exp <= 22'd2696823;
                12'd1162: exp <= 22'd2695657;
                12'd1163: exp <= 22'd2694491;
                12'd1164: exp <= 22'd2693326;
                12'd1165: exp <= 22'd2692160;
                12'd1166: exp <= 22'd2690995;
                12'd1167: exp <= 22'd2689830;
                12'd1168: exp <= 22'd2688665;
                12'd1169: exp <= 22'd2687500;
                12'd1170: exp <= 22'd2686336;
                12'd1171: exp <= 22'd2685172;
                12'd1172: exp <= 22'd2684008;
                12'd1173: exp <= 22'd2682844;
                12'd1174: exp <= 22'd2681680;
                12'd1175: exp <= 22'd2680517;
                12'd1176: exp <= 22'd2679353;
                12'd1177: exp <= 22'd2678190;
                12'd1178: exp <= 22'd2677027;
                12'd1179: exp <= 22'd2675865;
                12'd1180: exp <= 22'd2674702;
                12'd1181: exp <= 22'd2673540;
                12'd1182: exp <= 22'd2672378;
                12'd1183: exp <= 22'd2671216;
                12'd1184: exp <= 22'd2670054;
                12'd1185: exp <= 22'd2668892;
                12'd1186: exp <= 22'd2667731;
                12'd1187: exp <= 22'd2666570;
                12'd1188: exp <= 22'd2665409;
                12'd1189: exp <= 22'd2664248;
                12'd1190: exp <= 22'd2663088;
                12'd1191: exp <= 22'd2661927;
                12'd1192: exp <= 22'd2660767;
                12'd1193: exp <= 22'd2659607;
                12'd1194: exp <= 22'd2658448;
                12'd1195: exp <= 22'd2657288;
                12'd1196: exp <= 22'd2656129;
                12'd1197: exp <= 22'd2654969;
                12'd1198: exp <= 22'd2653810;
                12'd1199: exp <= 22'd2652652;
                12'd1200: exp <= 22'd2651493;
                12'd1201: exp <= 22'd2650335;
                12'd1202: exp <= 22'd2649177;
                12'd1203: exp <= 22'd2648019;
                12'd1204: exp <= 22'd2646861;
                12'd1205: exp <= 22'd2645703;
                12'd1206: exp <= 22'd2644546;
                12'd1207: exp <= 22'd2643389;
                12'd1208: exp <= 22'd2642232;
                12'd1209: exp <= 22'd2641075;
                12'd1210: exp <= 22'd2639918;
                12'd1211: exp <= 22'd2638762;
                12'd1212: exp <= 22'd2637605;
                12'd1213: exp <= 22'd2636449;
                12'd1214: exp <= 22'd2635294;
                12'd1215: exp <= 22'd2634138;
                12'd1216: exp <= 22'd2632982;
                12'd1217: exp <= 22'd2631827;
                12'd1218: exp <= 22'd2630672;
                12'd1219: exp <= 22'd2629517;
                12'd1220: exp <= 22'd2628363;
                12'd1221: exp <= 22'd2627208;
                12'd1222: exp <= 22'd2626054;
                12'd1223: exp <= 22'd2624900;
                12'd1224: exp <= 22'd2623746;
                12'd1225: exp <= 22'd2622592;
                12'd1226: exp <= 22'd2621439;
                12'd1227: exp <= 22'd2620285;
                12'd1228: exp <= 22'd2619132;
                12'd1229: exp <= 22'd2617979;
                12'd1230: exp <= 22'd2616827;
                12'd1231: exp <= 22'd2615674;
                12'd1232: exp <= 22'd2614522;
                12'd1233: exp <= 22'd2613370;
                12'd1234: exp <= 22'd2612218;
                12'd1235: exp <= 22'd2611066;
                12'd1236: exp <= 22'd2609915;
                12'd1237: exp <= 22'd2608763;
                12'd1238: exp <= 22'd2607612;
                12'd1239: exp <= 22'd2606461;
                12'd1240: exp <= 22'd2605310;
                12'd1241: exp <= 22'd2604160;
                12'd1242: exp <= 22'd2603009;
                12'd1243: exp <= 22'd2601859;
                12'd1244: exp <= 22'd2600709;
                12'd1245: exp <= 22'd2599559;
                12'd1246: exp <= 22'd2598410;
                12'd1247: exp <= 22'd2597260;
                12'd1248: exp <= 22'd2596111;
                12'd1249: exp <= 22'd2594962;
                12'd1250: exp <= 22'd2593813;
                12'd1251: exp <= 22'd2592665;
                12'd1252: exp <= 22'd2591516;
                12'd1253: exp <= 22'd2590368;
                12'd1254: exp <= 22'd2589220;
                12'd1255: exp <= 22'd2588072;
                12'd1256: exp <= 22'd2586925;
                12'd1257: exp <= 22'd2585777;
                12'd1258: exp <= 22'd2584630;
                12'd1259: exp <= 22'd2583483;
                12'd1260: exp <= 22'd2582336;
                12'd1261: exp <= 22'd2581189;
                12'd1262: exp <= 22'd2580043;
                12'd1263: exp <= 22'd2578896;
                12'd1264: exp <= 22'd2577750;
                12'd1265: exp <= 22'd2576604;
                12'd1266: exp <= 22'd2575459;
                12'd1267: exp <= 22'd2574313;
                12'd1268: exp <= 22'd2573168;
                12'd1269: exp <= 22'd2572023;
                12'd1270: exp <= 22'd2570878;
                12'd1271: exp <= 22'd2569733;
                12'd1272: exp <= 22'd2568588;
                12'd1273: exp <= 22'd2567444;
                12'd1274: exp <= 22'd2566300;
                12'd1275: exp <= 22'd2565156;
                12'd1276: exp <= 22'd2564012;
                12'd1277: exp <= 22'd2562869;
                12'd1278: exp <= 22'd2561725;
                12'd1279: exp <= 22'd2560582;
                12'd1280: exp <= 22'd2559439;
                12'd1281: exp <= 22'd2558296;
                12'd1282: exp <= 22'd2557154;
                12'd1283: exp <= 22'd2556011;
                12'd1284: exp <= 22'd2554869;
                12'd1285: exp <= 22'd2553727;
                12'd1286: exp <= 22'd2552585;
                12'd1287: exp <= 22'd2551443;
                12'd1288: exp <= 22'd2550302;
                12'd1289: exp <= 22'd2549161;
                12'd1290: exp <= 22'd2548020;
                12'd1291: exp <= 22'd2546879;
                12'd1292: exp <= 22'd2545738;
                12'd1293: exp <= 22'd2544598;
                12'd1294: exp <= 22'd2543457;
                12'd1295: exp <= 22'd2542317;
                12'd1296: exp <= 22'd2541177;
                12'd1297: exp <= 22'd2540038;
                12'd1298: exp <= 22'd2538898;
                12'd1299: exp <= 22'd2537759;
                12'd1300: exp <= 22'd2536620;
                12'd1301: exp <= 22'd2535481;
                12'd1302: exp <= 22'd2534342;
                12'd1303: exp <= 22'd2533203;
                12'd1304: exp <= 22'd2532065;
                12'd1305: exp <= 22'd2530927;
                12'd1306: exp <= 22'd2529789;
                12'd1307: exp <= 22'd2528651;
                12'd1308: exp <= 22'd2527513;
                12'd1309: exp <= 22'd2526376;
                12'd1310: exp <= 22'd2525239;
                12'd1311: exp <= 22'd2524102;
                12'd1312: exp <= 22'd2522965;
                12'd1313: exp <= 22'd2521828;
                12'd1314: exp <= 22'd2520692;
                12'd1315: exp <= 22'd2519556;
                12'd1316: exp <= 22'd2518420;
                12'd1317: exp <= 22'd2517284;
                12'd1318: exp <= 22'd2516148;
                12'd1319: exp <= 22'd2515013;
                12'd1320: exp <= 22'd2513877;
                12'd1321: exp <= 22'd2512742;
                12'd1322: exp <= 22'd2511607;
                12'd1323: exp <= 22'd2510473;
                12'd1324: exp <= 22'd2509338;
                12'd1325: exp <= 22'd2508204;
                12'd1326: exp <= 22'd2507070;
                12'd1327: exp <= 22'd2505936;
                12'd1328: exp <= 22'd2504802;
                12'd1329: exp <= 22'd2503668;
                12'd1330: exp <= 22'd2502535;
                12'd1331: exp <= 22'd2501402;
                12'd1332: exp <= 22'd2500269;
                12'd1333: exp <= 22'd2499136;
                12'd1334: exp <= 22'd2498003;
                12'd1335: exp <= 22'd2496871;
                12'd1336: exp <= 22'd2495739;
                12'd1337: exp <= 22'd2494607;
                12'd1338: exp <= 22'd2493475;
                12'd1339: exp <= 22'd2492343;
                12'd1340: exp <= 22'd2491212;
                12'd1341: exp <= 22'd2490080;
                12'd1342: exp <= 22'd2488949;
                12'd1343: exp <= 22'd2487818;
                12'd1344: exp <= 22'd2486688;
                12'd1345: exp <= 22'd2485557;
                12'd1346: exp <= 22'd2484427;
                12'd1347: exp <= 22'd2483297;
                12'd1348: exp <= 22'd2482167;
                12'd1349: exp <= 22'd2481037;
                12'd1350: exp <= 22'd2479908;
                12'd1351: exp <= 22'd2478778;
                12'd1352: exp <= 22'd2477649;
                12'd1353: exp <= 22'd2476520;
                12'd1354: exp <= 22'd2475391;
                12'd1355: exp <= 22'd2474263;
                12'd1356: exp <= 22'd2473134;
                12'd1357: exp <= 22'd2472006;
                12'd1358: exp <= 22'd2470878;
                12'd1359: exp <= 22'd2469750;
                12'd1360: exp <= 22'd2468623;
                12'd1361: exp <= 22'd2467495;
                12'd1362: exp <= 22'd2466368;
                12'd1363: exp <= 22'd2465241;
                12'd1364: exp <= 22'd2464114;
                12'd1365: exp <= 22'd2462987;
                12'd1366: exp <= 22'd2461861;
                12'd1367: exp <= 22'd2460735;
                12'd1368: exp <= 22'd2459609;
                12'd1369: exp <= 22'd2458483;
                12'd1370: exp <= 22'd2457357;
                12'd1371: exp <= 22'd2456231;
                12'd1372: exp <= 22'd2455106;
                12'd1373: exp <= 22'd2453981;
                12'd1374: exp <= 22'd2452856;
                12'd1375: exp <= 22'd2451731;
                12'd1376: exp <= 22'd2450607;
                12'd1377: exp <= 22'd2449482;
                12'd1378: exp <= 22'd2448358;
                12'd1379: exp <= 22'd2447234;
                12'd1380: exp <= 22'd2446110;
                12'd1381: exp <= 22'd2444987;
                12'd1382: exp <= 22'd2443863;
                12'd1383: exp <= 22'd2442740;
                12'd1384: exp <= 22'd2441617;
                12'd1385: exp <= 22'd2440494;
                12'd1386: exp <= 22'd2439371;
                12'd1387: exp <= 22'd2438249;
                12'd1388: exp <= 22'd2437126;
                12'd1389: exp <= 22'd2436004;
                12'd1390: exp <= 22'd2434882;
                12'd1391: exp <= 22'd2433761;
                12'd1392: exp <= 22'd2432639;
                12'd1393: exp <= 22'd2431518;
                12'd1394: exp <= 22'd2430397;
                12'd1395: exp <= 22'd2429276;
                12'd1396: exp <= 22'd2428155;
                12'd1397: exp <= 22'd2427034;
                12'd1398: exp <= 22'd2425914;
                12'd1399: exp <= 22'd2424794;
                12'd1400: exp <= 22'd2423674;
                12'd1401: exp <= 22'd2422554;
                12'd1402: exp <= 22'd2421434;
                12'd1403: exp <= 22'd2420315;
                12'd1404: exp <= 22'd2419195;
                12'd1405: exp <= 22'd2418076;
                12'd1406: exp <= 22'd2416957;
                12'd1407: exp <= 22'd2415839;
                12'd1408: exp <= 22'd2414720;
                12'd1409: exp <= 22'd2413602;
                12'd1410: exp <= 22'd2412484;
                12'd1411: exp <= 22'd2411366;
                12'd1412: exp <= 22'd2410248;
                12'd1413: exp <= 22'd2409131;
                12'd1414: exp <= 22'd2408013;
                12'd1415: exp <= 22'd2406896;
                12'd1416: exp <= 22'd2405779;
                12'd1417: exp <= 22'd2404662;
                12'd1418: exp <= 22'd2403546;
                12'd1419: exp <= 22'd2402429;
                12'd1420: exp <= 22'd2401313;
                12'd1421: exp <= 22'd2400197;
                12'd1422: exp <= 22'd2399081;
                12'd1423: exp <= 22'd2397965;
                12'd1424: exp <= 22'd2396850;
                12'd1425: exp <= 22'd2395735;
                12'd1426: exp <= 22'd2394619;
                12'd1427: exp <= 22'd2393504;
                12'd1428: exp <= 22'd2392390;
                12'd1429: exp <= 22'd2391275;
                12'd1430: exp <= 22'd2390161;
                12'd1431: exp <= 22'd2389047;
                12'd1432: exp <= 22'd2387933;
                12'd1433: exp <= 22'd2386819;
                12'd1434: exp <= 22'd2385705;
                12'd1435: exp <= 22'd2384592;
                12'd1436: exp <= 22'd2383479;
                12'd1437: exp <= 22'd2382366;
                12'd1438: exp <= 22'd2381253;
                12'd1439: exp <= 22'd2380140;
                12'd1440: exp <= 22'd2379028;
                12'd1441: exp <= 22'd2377915;
                12'd1442: exp <= 22'd2376803;
                12'd1443: exp <= 22'd2375691;
                12'd1444: exp <= 22'd2374580;
                12'd1445: exp <= 22'd2373468;
                12'd1446: exp <= 22'd2372357;
                12'd1447: exp <= 22'd2371246;
                12'd1448: exp <= 22'd2370135;
                12'd1449: exp <= 22'd2369024;
                12'd1450: exp <= 22'd2367913;
                12'd1451: exp <= 22'd2366803;
                12'd1452: exp <= 22'd2365693;
                12'd1453: exp <= 22'd2364583;
                12'd1454: exp <= 22'd2363473;
                12'd1455: exp <= 22'd2362363;
                12'd1456: exp <= 22'd2361254;
                12'd1457: exp <= 22'd2360145;
                12'd1458: exp <= 22'd2359035;
                12'd1459: exp <= 22'd2357927;
                12'd1460: exp <= 22'd2356818;
                12'd1461: exp <= 22'd2355709;
                12'd1462: exp <= 22'd2354601;
                12'd1463: exp <= 22'd2353493;
                12'd1464: exp <= 22'd2352385;
                12'd1465: exp <= 22'd2351277;
                12'd1466: exp <= 22'd2350170;
                12'd1467: exp <= 22'd2349062;
                12'd1468: exp <= 22'd2347955;
                12'd1469: exp <= 22'd2346848;
                12'd1470: exp <= 22'd2345741;
                12'd1471: exp <= 22'd2344634;
                12'd1472: exp <= 22'd2343528;
                12'd1473: exp <= 22'd2342422;
                12'd1474: exp <= 22'd2341316;
                12'd1475: exp <= 22'd2340210;
                12'd1476: exp <= 22'd2339104;
                12'd1477: exp <= 22'd2337998;
                12'd1478: exp <= 22'd2336893;
                12'd1479: exp <= 22'd2335788;
                12'd1480: exp <= 22'd2334683;
                12'd1481: exp <= 22'd2333578;
                12'd1482: exp <= 22'd2332474;
                12'd1483: exp <= 22'd2331369;
                12'd1484: exp <= 22'd2330265;
                12'd1485: exp <= 22'd2329161;
                12'd1486: exp <= 22'd2328057;
                12'd1487: exp <= 22'd2326953;
                12'd1488: exp <= 22'd2325850;
                12'd1489: exp <= 22'd2324747;
                12'd1490: exp <= 22'd2323644;
                12'd1491: exp <= 22'd2322541;
                12'd1492: exp <= 22'd2321438;
                12'd1493: exp <= 22'd2320335;
                12'd1494: exp <= 22'd2319233;
                12'd1495: exp <= 22'd2318131;
                12'd1496: exp <= 22'd2317029;
                12'd1497: exp <= 22'd2315927;
                12'd1498: exp <= 22'd2314826;
                12'd1499: exp <= 22'd2313724;
                12'd1500: exp <= 22'd2312623;
                12'd1501: exp <= 22'd2311522;
                12'd1502: exp <= 22'd2310421;
                12'd1503: exp <= 22'd2309320;
                12'd1504: exp <= 22'd2308220;
                12'd1505: exp <= 22'd2307120;
                12'd1506: exp <= 22'd2306019;
                12'd1507: exp <= 22'd2304920;
                12'd1508: exp <= 22'd2303820;
                12'd1509: exp <= 22'd2302720;
                12'd1510: exp <= 22'd2301621;
                12'd1511: exp <= 22'd2300522;
                12'd1512: exp <= 22'd2299423;
                12'd1513: exp <= 22'd2298324;
                12'd1514: exp <= 22'd2297225;
                12'd1515: exp <= 22'd2296127;
                12'd1516: exp <= 22'd2295029;
                12'd1517: exp <= 22'd2293930;
                12'd1518: exp <= 22'd2292833;
                12'd1519: exp <= 22'd2291735;
                12'd1520: exp <= 22'd2290637;
                12'd1521: exp <= 22'd2289540;
                12'd1522: exp <= 22'd2288443;
                12'd1523: exp <= 22'd2287346;
                12'd1524: exp <= 22'd2286249;
                12'd1525: exp <= 22'd2285153;
                12'd1526: exp <= 22'd2284056;
                12'd1527: exp <= 22'd2282960;
                12'd1528: exp <= 22'd2281864;
                12'd1529: exp <= 22'd2280768;
                12'd1530: exp <= 22'd2279673;
                12'd1531: exp <= 22'd2278577;
                12'd1532: exp <= 22'd2277482;
                12'd1533: exp <= 22'd2276387;
                12'd1534: exp <= 22'd2275292;
                12'd1535: exp <= 22'd2274197;
                12'd1536: exp <= 22'd2273102;
                12'd1537: exp <= 22'd2272008;
                12'd1538: exp <= 22'd2270914;
                12'd1539: exp <= 22'd2269820;
                12'd1540: exp <= 22'd2268726;
                12'd1541: exp <= 22'd2267633;
                12'd1542: exp <= 22'd2266539;
                12'd1543: exp <= 22'd2265446;
                12'd1544: exp <= 22'd2264353;
                12'd1545: exp <= 22'd2263260;
                12'd1546: exp <= 22'd2262167;
                12'd1547: exp <= 22'd2261075;
                12'd1548: exp <= 22'd2259982;
                12'd1549: exp <= 22'd2258890;
                12'd1550: exp <= 22'd2257798;
                12'd1551: exp <= 22'd2256707;
                12'd1552: exp <= 22'd2255615;
                12'd1553: exp <= 22'd2254524;
                12'd1554: exp <= 22'd2253432;
                12'd1555: exp <= 22'd2252341;
                12'd1556: exp <= 22'd2251251;
                12'd1557: exp <= 22'd2250160;
                12'd1558: exp <= 22'd2249069;
                12'd1559: exp <= 22'd2247979;
                12'd1560: exp <= 22'd2246889;
                12'd1561: exp <= 22'd2245799;
                12'd1562: exp <= 22'd2244709;
                12'd1563: exp <= 22'd2243620;
                12'd1564: exp <= 22'd2242530;
                12'd1565: exp <= 22'd2241441;
                12'd1566: exp <= 22'd2240352;
                12'd1567: exp <= 22'd2239263;
                12'd1568: exp <= 22'd2238175;
                12'd1569: exp <= 22'd2237086;
                12'd1570: exp <= 22'd2235998;
                12'd1571: exp <= 22'd2234910;
                12'd1572: exp <= 22'd2233822;
                12'd1573: exp <= 22'd2232734;
                12'd1574: exp <= 22'd2231647;
                12'd1575: exp <= 22'd2230560;
                12'd1576: exp <= 22'd2229472;
                12'd1577: exp <= 22'd2228385;
                12'd1578: exp <= 22'd2227299;
                12'd1579: exp <= 22'd2226212;
                12'd1580: exp <= 22'd2225126;
                12'd1581: exp <= 22'd2224039;
                12'd1582: exp <= 22'd2222953;
                12'd1583: exp <= 22'd2221867;
                12'd1584: exp <= 22'd2220782;
                12'd1585: exp <= 22'd2219696;
                12'd1586: exp <= 22'd2218611;
                12'd1587: exp <= 22'd2217526;
                12'd1588: exp <= 22'd2216441;
                12'd1589: exp <= 22'd2215356;
                12'd1590: exp <= 22'd2214271;
                12'd1591: exp <= 22'd2213187;
                12'd1592: exp <= 22'd2212103;
                12'd1593: exp <= 22'd2211019;
                12'd1594: exp <= 22'd2209935;
                12'd1595: exp <= 22'd2208851;
                12'd1596: exp <= 22'd2207768;
                12'd1597: exp <= 22'd2206684;
                12'd1598: exp <= 22'd2205601;
                12'd1599: exp <= 22'd2204518;
                12'd1600: exp <= 22'd2203436;
                12'd1601: exp <= 22'd2202353;
                12'd1602: exp <= 22'd2201271;
                12'd1603: exp <= 22'd2200189;
                12'd1604: exp <= 22'd2199107;
                12'd1605: exp <= 22'd2198025;
                12'd1606: exp <= 22'd2196943;
                12'd1607: exp <= 22'd2195862;
                12'd1608: exp <= 22'd2194780;
                12'd1609: exp <= 22'd2193699;
                12'd1610: exp <= 22'd2192618;
                12'd1611: exp <= 22'd2191537;
                12'd1612: exp <= 22'd2190457;
                12'd1613: exp <= 22'd2189377;
                12'd1614: exp <= 22'd2188296;
                12'd1615: exp <= 22'd2187216;
                12'd1616: exp <= 22'd2186137;
                12'd1617: exp <= 22'd2185057;
                12'd1618: exp <= 22'd2183977;
                12'd1619: exp <= 22'd2182898;
                12'd1620: exp <= 22'd2181819;
                12'd1621: exp <= 22'd2180740;
                12'd1622: exp <= 22'd2179661;
                12'd1623: exp <= 22'd2178583;
                12'd1624: exp <= 22'd2177505;
                12'd1625: exp <= 22'd2176426;
                12'd1626: exp <= 22'd2175348;
                12'd1627: exp <= 22'd2174271;
                12'd1628: exp <= 22'd2173193;
                12'd1629: exp <= 22'd2172115;
                12'd1630: exp <= 22'd2171038;
                12'd1631: exp <= 22'd2169961;
                12'd1632: exp <= 22'd2168884;
                12'd1633: exp <= 22'd2167807;
                12'd1634: exp <= 22'd2166731;
                12'd1635: exp <= 22'd2165655;
                12'd1636: exp <= 22'd2164578;
                12'd1637: exp <= 22'd2163502;
                12'd1638: exp <= 22'd2162427;
                12'd1639: exp <= 22'd2161351;
                12'd1640: exp <= 22'd2160276;
                12'd1641: exp <= 22'd2159200;
                12'd1642: exp <= 22'd2158125;
                12'd1643: exp <= 22'd2157050;
                12'd1644: exp <= 22'd2155976;
                12'd1645: exp <= 22'd2154901;
                12'd1646: exp <= 22'd2153827;
                12'd1647: exp <= 22'd2152752;
                12'd1648: exp <= 22'd2151678;
                12'd1649: exp <= 22'd2150605;
                12'd1650: exp <= 22'd2149531;
                12'd1651: exp <= 22'd2148458;
                12'd1652: exp <= 22'd2147384;
                12'd1653: exp <= 22'd2146311;
                12'd1654: exp <= 22'd2145238;
                12'd1655: exp <= 22'd2144166;
                12'd1656: exp <= 22'd2143093;
                12'd1657: exp <= 22'd2142021;
                12'd1658: exp <= 22'd2140949;
                12'd1659: exp <= 22'd2139877;
                12'd1660: exp <= 22'd2138805;
                12'd1661: exp <= 22'd2137733;
                12'd1662: exp <= 22'd2136662;
                12'd1663: exp <= 22'd2135590;
                12'd1664: exp <= 22'd2134519;
                12'd1665: exp <= 22'd2133448;
                12'd1666: exp <= 22'd2132378;
                12'd1667: exp <= 22'd2131307;
                12'd1668: exp <= 22'd2130237;
                12'd1669: exp <= 22'd2129167;
                12'd1670: exp <= 22'd2128097;
                12'd1671: exp <= 22'd2127027;
                12'd1672: exp <= 22'd2125957;
                12'd1673: exp <= 22'd2124888;
                12'd1674: exp <= 22'd2123818;
                12'd1675: exp <= 22'd2122749;
                12'd1676: exp <= 22'd2121680;
                12'd1677: exp <= 22'd2120612;
                12'd1678: exp <= 22'd2119543;
                12'd1679: exp <= 22'd2118475;
                12'd1680: exp <= 22'd2117407;
                12'd1681: exp <= 22'd2116339;
                12'd1682: exp <= 22'd2115271;
                12'd1683: exp <= 22'd2114203;
                12'd1684: exp <= 22'd2113136;
                12'd1685: exp <= 22'd2112068;
                12'd1686: exp <= 22'd2111001;
                12'd1687: exp <= 22'd2109934;
                12'd1688: exp <= 22'd2108867;
                12'd1689: exp <= 22'd2107801;
                12'd1690: exp <= 22'd2106735;
                12'd1691: exp <= 22'd2105668;
                12'd1692: exp <= 22'd2104602;
                12'd1693: exp <= 22'd2103536;
                12'd1694: exp <= 22'd2102471;
                12'd1695: exp <= 22'd2101405;
                12'd1696: exp <= 22'd2100340;
                12'd1697: exp <= 22'd2099275;
                12'd1698: exp <= 22'd2098210;
                12'd1699: exp <= 22'd2097145;
                12'd1700: exp <= 22'd2096081;
                12'd1701: exp <= 22'd2095016;
                12'd1702: exp <= 22'd2093952;
                12'd1703: exp <= 22'd2092888;
                12'd1704: exp <= 22'd2091824;
                12'd1705: exp <= 22'd2090760;
                12'd1706: exp <= 22'd2089697;
                12'd1707: exp <= 22'd2088634;
                12'd1708: exp <= 22'd2087570;
                12'd1709: exp <= 22'd2086507;
                12'd1710: exp <= 22'd2085445;
                12'd1711: exp <= 22'd2084382;
                12'd1712: exp <= 22'd2083320;
                12'd1713: exp <= 22'd2082257;
                12'd1714: exp <= 22'd2081195;
                12'd1715: exp <= 22'd2080133;
                12'd1716: exp <= 22'd2079072;
                12'd1717: exp <= 22'd2078010;
                12'd1718: exp <= 22'd2076949;
                12'd1719: exp <= 22'd2075888;
                12'd1720: exp <= 22'd2074827;
                12'd1721: exp <= 22'd2073766;
                12'd1722: exp <= 22'd2072705;
                12'd1723: exp <= 22'd2071645;
                12'd1724: exp <= 22'd2070585;
                12'd1725: exp <= 22'd2069524;
                12'd1726: exp <= 22'd2068465;
                12'd1727: exp <= 22'd2067405;
                12'd1728: exp <= 22'd2066345;
                12'd1729: exp <= 22'd2065286;
                12'd1730: exp <= 22'd2064227;
                12'd1731: exp <= 22'd2063168;
                12'd1732: exp <= 22'd2062109;
                12'd1733: exp <= 22'd2061050;
                12'd1734: exp <= 22'd2059992;
                12'd1735: exp <= 22'd2058933;
                12'd1736: exp <= 22'd2057875;
                12'd1737: exp <= 22'd2056817;
                12'd1738: exp <= 22'd2055760;
                12'd1739: exp <= 22'd2054702;
                12'd1740: exp <= 22'd2053645;
                12'd1741: exp <= 22'd2052587;
                12'd1742: exp <= 22'd2051530;
                12'd1743: exp <= 22'd2050474;
                12'd1744: exp <= 22'd2049417;
                12'd1745: exp <= 22'd2048360;
                12'd1746: exp <= 22'd2047304;
                12'd1747: exp <= 22'd2046248;
                12'd1748: exp <= 22'd2045192;
                12'd1749: exp <= 22'd2044136;
                12'd1750: exp <= 22'd2043081;
                12'd1751: exp <= 22'd2042025;
                12'd1752: exp <= 22'd2040970;
                12'd1753: exp <= 22'd2039915;
                12'd1754: exp <= 22'd2038860;
                12'd1755: exp <= 22'd2037805;
                12'd1756: exp <= 22'd2036751;
                12'd1757: exp <= 22'd2035696;
                12'd1758: exp <= 22'd2034642;
                12'd1759: exp <= 22'd2033588;
                12'd1760: exp <= 22'd2032534;
                12'd1761: exp <= 22'd2031481;
                12'd1762: exp <= 22'd2030427;
                12'd1763: exp <= 22'd2029374;
                12'd1764: exp <= 22'd2028321;
                12'd1765: exp <= 22'd2027268;
                12'd1766: exp <= 22'd2026215;
                12'd1767: exp <= 22'd2025162;
                12'd1768: exp <= 22'd2024110;
                12'd1769: exp <= 22'd2023058;
                12'd1770: exp <= 22'd2022006;
                12'd1771: exp <= 22'd2020954;
                12'd1772: exp <= 22'd2019902;
                12'd1773: exp <= 22'd2018851;
                12'd1774: exp <= 22'd2017799;
                12'd1775: exp <= 22'd2016748;
                12'd1776: exp <= 22'd2015697;
                12'd1777: exp <= 22'd2014646;
                12'd1778: exp <= 22'd2013596;
                12'd1779: exp <= 22'd2012545;
                12'd1780: exp <= 22'd2011495;
                12'd1781: exp <= 22'd2010445;
                12'd1782: exp <= 22'd2009395;
                12'd1783: exp <= 22'd2008345;
                12'd1784: exp <= 22'd2007296;
                12'd1785: exp <= 22'd2006246;
                12'd1786: exp <= 22'd2005197;
                12'd1787: exp <= 22'd2004148;
                12'd1788: exp <= 22'd2003099;
                12'd1789: exp <= 22'd2002051;
                12'd1790: exp <= 22'd2001002;
                12'd1791: exp <= 22'd1999954;
                12'd1792: exp <= 22'd1998906;
                12'd1793: exp <= 22'd1997858;
                12'd1794: exp <= 22'd1996810;
                12'd1795: exp <= 22'd1995762;
                12'd1796: exp <= 22'd1994715;
                12'd1797: exp <= 22'd1993668;
                12'd1798: exp <= 22'd1992621;
                12'd1799: exp <= 22'd1991574;
                12'd1800: exp <= 22'd1990527;
                12'd1801: exp <= 22'd1989480;
                12'd1802: exp <= 22'd1988434;
                12'd1803: exp <= 22'd1987388;
                12'd1804: exp <= 22'd1986342;
                12'd1805: exp <= 22'd1985296;
                12'd1806: exp <= 22'd1984250;
                12'd1807: exp <= 22'd1983205;
                12'd1808: exp <= 22'd1982160;
                12'd1809: exp <= 22'd1981114;
                12'd1810: exp <= 22'd1980070;
                12'd1811: exp <= 22'd1979025;
                12'd1812: exp <= 22'd1977980;
                12'd1813: exp <= 22'd1976936;
                12'd1814: exp <= 22'd1975891;
                12'd1815: exp <= 22'd1974847;
                12'd1816: exp <= 22'd1973804;
                12'd1817: exp <= 22'd1972760;
                12'd1818: exp <= 22'd1971716;
                12'd1819: exp <= 22'd1970673;
                12'd1820: exp <= 22'd1969630;
                12'd1821: exp <= 22'd1968587;
                12'd1822: exp <= 22'd1967544;
                12'd1823: exp <= 22'd1966501;
                12'd1824: exp <= 22'd1965459;
                12'd1825: exp <= 22'd1964416;
                12'd1826: exp <= 22'd1963374;
                12'd1827: exp <= 22'd1962332;
                12'd1828: exp <= 22'd1961291;
                12'd1829: exp <= 22'd1960249;
                12'd1830: exp <= 22'd1959208;
                12'd1831: exp <= 22'd1958166;
                12'd1832: exp <= 22'd1957125;
                12'd1833: exp <= 22'd1956084;
                12'd1834: exp <= 22'd1955044;
                12'd1835: exp <= 22'd1954003;
                12'd1836: exp <= 22'd1952963;
                12'd1837: exp <= 22'd1951923;
                12'd1838: exp <= 22'd1950883;
                12'd1839: exp <= 22'd1949843;
                12'd1840: exp <= 22'd1948803;
                12'd1841: exp <= 22'd1947764;
                12'd1842: exp <= 22'd1946724;
                12'd1843: exp <= 22'd1945685;
                12'd1844: exp <= 22'd1944646;
                12'd1845: exp <= 22'd1943607;
                12'd1846: exp <= 22'd1942569;
                12'd1847: exp <= 22'd1941530;
                12'd1848: exp <= 22'd1940492;
                12'd1849: exp <= 22'd1939454;
                12'd1850: exp <= 22'd1938416;
                12'd1851: exp <= 22'd1937378;
                12'd1852: exp <= 22'd1936341;
                12'd1853: exp <= 22'd1935304;
                12'd1854: exp <= 22'd1934266;
                12'd1855: exp <= 22'd1933229;
                12'd1856: exp <= 22'd1932193;
                12'd1857: exp <= 22'd1931156;
                12'd1858: exp <= 22'd1930119;
                12'd1859: exp <= 22'd1929083;
                12'd1860: exp <= 22'd1928047;
                12'd1861: exp <= 22'd1927011;
                12'd1862: exp <= 22'd1925975;
                12'd1863: exp <= 22'd1924939;
                12'd1864: exp <= 22'd1923904;
                12'd1865: exp <= 22'd1922869;
                12'd1866: exp <= 22'd1921834;
                12'd1867: exp <= 22'd1920799;
                12'd1868: exp <= 22'd1919764;
                12'd1869: exp <= 22'd1918729;
                12'd1870: exp <= 22'd1917695;
                12'd1871: exp <= 22'd1916661;
                12'd1872: exp <= 22'd1915627;
                12'd1873: exp <= 22'd1914593;
                12'd1874: exp <= 22'd1913559;
                12'd1875: exp <= 22'd1912526;
                12'd1876: exp <= 22'd1911492;
                12'd1877: exp <= 22'd1910459;
                12'd1878: exp <= 22'd1909426;
                12'd1879: exp <= 22'd1908393;
                12'd1880: exp <= 22'd1907361;
                12'd1881: exp <= 22'd1906328;
                12'd1882: exp <= 22'd1905296;
                12'd1883: exp <= 22'd1904264;
                12'd1884: exp <= 22'd1903232;
                12'd1885: exp <= 22'd1902200;
                12'd1886: exp <= 22'd1901169;
                12'd1887: exp <= 22'd1900137;
                12'd1888: exp <= 22'd1899106;
                12'd1889: exp <= 22'd1898075;
                12'd1890: exp <= 22'd1897044;
                12'd1891: exp <= 22'd1896013;
                12'd1892: exp <= 22'd1894983;
                12'd1893: exp <= 22'd1893952;
                12'd1894: exp <= 22'd1892922;
                12'd1895: exp <= 22'd1891892;
                12'd1896: exp <= 22'd1890862;
                12'd1897: exp <= 22'd1889833;
                12'd1898: exp <= 22'd1888803;
                12'd1899: exp <= 22'd1887774;
                12'd1900: exp <= 22'd1886745;
                12'd1901: exp <= 22'd1885716;
                12'd1902: exp <= 22'd1884687;
                12'd1903: exp <= 22'd1883658;
                12'd1904: exp <= 22'd1882630;
                12'd1905: exp <= 22'd1881601;
                12'd1906: exp <= 22'd1880573;
                12'd1907: exp <= 22'd1879545;
                12'd1908: exp <= 22'd1878518;
                12'd1909: exp <= 22'd1877490;
                12'd1910: exp <= 22'd1876463;
                12'd1911: exp <= 22'd1875435;
                12'd1912: exp <= 22'd1874408;
                12'd1913: exp <= 22'd1873381;
                12'd1914: exp <= 22'd1872355;
                12'd1915: exp <= 22'd1871328;
                12'd1916: exp <= 22'd1870302;
                12'd1917: exp <= 22'd1869276;
                12'd1918: exp <= 22'd1868249;
                12'd1919: exp <= 22'd1867224;
                12'd1920: exp <= 22'd1866198;
                12'd1921: exp <= 22'd1865172;
                12'd1922: exp <= 22'd1864147;
                12'd1923: exp <= 22'd1863122;
                12'd1924: exp <= 22'd1862097;
                12'd1925: exp <= 22'd1861072;
                12'd1926: exp <= 22'd1860048;
                12'd1927: exp <= 22'd1859023;
                12'd1928: exp <= 22'd1857999;
                12'd1929: exp <= 22'd1856975;
                12'd1930: exp <= 22'd1855951;
                12'd1931: exp <= 22'd1854927;
                12'd1932: exp <= 22'd1853903;
                12'd1933: exp <= 22'd1852880;
                12'd1934: exp <= 22'd1851857;
                12'd1935: exp <= 22'd1850834;
                12'd1936: exp <= 22'd1849811;
                12'd1937: exp <= 22'd1848788;
                12'd1938: exp <= 22'd1847765;
                12'd1939: exp <= 22'd1846743;
                12'd1940: exp <= 22'd1845721;
                12'd1941: exp <= 22'd1844699;
                12'd1942: exp <= 22'd1843677;
                12'd1943: exp <= 22'd1842655;
                12'd1944: exp <= 22'd1841634;
                12'd1945: exp <= 22'd1840612;
                12'd1946: exp <= 22'd1839591;
                12'd1947: exp <= 22'd1838570;
                12'd1948: exp <= 22'd1837549;
                12'd1949: exp <= 22'd1836529;
                12'd1950: exp <= 22'd1835508;
                12'd1951: exp <= 22'd1834488;
                12'd1952: exp <= 22'd1833468;
                12'd1953: exp <= 22'd1832448;
                12'd1954: exp <= 22'd1831428;
                12'd1955: exp <= 22'd1830408;
                12'd1956: exp <= 22'd1829389;
                12'd1957: exp <= 22'd1828370;
                12'd1958: exp <= 22'd1827351;
                12'd1959: exp <= 22'd1826332;
                12'd1960: exp <= 22'd1825313;
                12'd1961: exp <= 22'd1824294;
                12'd1962: exp <= 22'd1823276;
                12'd1963: exp <= 22'd1822258;
                12'd1964: exp <= 22'd1821240;
                12'd1965: exp <= 22'd1820222;
                12'd1966: exp <= 22'd1819204;
                12'd1967: exp <= 22'd1818186;
                12'd1968: exp <= 22'd1817169;
                12'd1969: exp <= 22'd1816152;
                12'd1970: exp <= 22'd1815135;
                12'd1971: exp <= 22'd1814118;
                12'd1972: exp <= 22'd1813101;
                12'd1973: exp <= 22'd1812085;
                12'd1974: exp <= 22'd1811068;
                12'd1975: exp <= 22'd1810052;
                12'd1976: exp <= 22'd1809036;
                12'd1977: exp <= 22'd1808020;
                12'd1978: exp <= 22'd1807005;
                12'd1979: exp <= 22'd1805989;
                12'd1980: exp <= 22'd1804974;
                12'd1981: exp <= 22'd1803959;
                12'd1982: exp <= 22'd1802944;
                12'd1983: exp <= 22'd1801929;
                12'd1984: exp <= 22'd1800914;
                12'd1985: exp <= 22'd1799900;
                12'd1986: exp <= 22'd1798886;
                12'd1987: exp <= 22'd1797871;
                12'd1988: exp <= 22'd1796858;
                12'd1989: exp <= 22'd1795844;
                12'd1990: exp <= 22'd1794830;
                12'd1991: exp <= 22'd1793817;
                12'd1992: exp <= 22'd1792803;
                12'd1993: exp <= 22'd1791790;
                12'd1994: exp <= 22'd1790777;
                12'd1995: exp <= 22'd1789765;
                12'd1996: exp <= 22'd1788752;
                12'd1997: exp <= 22'd1787740;
                12'd1998: exp <= 22'd1786728;
                12'd1999: exp <= 22'd1785715;
                12'd2000: exp <= 22'd1784704;
                12'd2001: exp <= 22'd1783692;
                12'd2002: exp <= 22'd1782680;
                12'd2003: exp <= 22'd1781669;
                12'd2004: exp <= 22'd1780658;
                12'd2005: exp <= 22'd1779647;
                12'd2006: exp <= 22'd1778636;
                12'd2007: exp <= 22'd1777625;
                12'd2008: exp <= 22'd1776615;
                12'd2009: exp <= 22'd1775604;
                12'd2010: exp <= 22'd1774594;
                12'd2011: exp <= 22'd1773584;
                12'd2012: exp <= 22'd1772574;
                12'd2013: exp <= 22'd1771565;
                12'd2014: exp <= 22'd1770555;
                12'd2015: exp <= 22'd1769546;
                12'd2016: exp <= 22'd1768537;
                12'd2017: exp <= 22'd1767528;
                12'd2018: exp <= 22'd1766519;
                12'd2019: exp <= 22'd1765510;
                12'd2020: exp <= 22'd1764502;
                12'd2021: exp <= 22'd1763493;
                12'd2022: exp <= 22'd1762485;
                12'd2023: exp <= 22'd1761477;
                12'd2024: exp <= 22'd1760470;
                12'd2025: exp <= 22'd1759462;
                12'd2026: exp <= 22'd1758455;
                12'd2027: exp <= 22'd1757447;
                12'd2028: exp <= 22'd1756440;
                12'd2029: exp <= 22'd1755433;
                12'd2030: exp <= 22'd1754427;
                12'd2031: exp <= 22'd1753420;
                12'd2032: exp <= 22'd1752413;
                12'd2033: exp <= 22'd1751407;
                12'd2034: exp <= 22'd1750401;
                12'd2035: exp <= 22'd1749395;
                12'd2036: exp <= 22'd1748390;
                12'd2037: exp <= 22'd1747384;
                12'd2038: exp <= 22'd1746379;
                12'd2039: exp <= 22'd1745373;
                12'd2040: exp <= 22'd1744368;
                12'd2041: exp <= 22'd1743363;
                12'd2042: exp <= 22'd1742359;
                12'd2043: exp <= 22'd1741354;
                12'd2044: exp <= 22'd1740350;
                12'd2045: exp <= 22'd1739346;
                12'd2046: exp <= 22'd1738341;
                12'd2047: exp <= 22'd1737338;
                12'd2048: exp <= 22'd1736334;
                12'd2049: exp <= 22'd1735330;
                12'd2050: exp <= 22'd1734327;
                12'd2051: exp <= 22'd1733324;
                12'd2052: exp <= 22'd1732321;
                12'd2053: exp <= 22'd1731318;
                12'd2054: exp <= 22'd1730315;
                12'd2055: exp <= 22'd1729313;
                12'd2056: exp <= 22'd1728310;
                12'd2057: exp <= 22'd1727308;
                12'd2058: exp <= 22'd1726306;
                12'd2059: exp <= 22'd1725304;
                12'd2060: exp <= 22'd1724303;
                12'd2061: exp <= 22'd1723301;
                12'd2062: exp <= 22'd1722300;
                12'd2063: exp <= 22'd1721299;
                12'd2064: exp <= 22'd1720298;
                12'd2065: exp <= 22'd1719297;
                12'd2066: exp <= 22'd1718296;
                12'd2067: exp <= 22'd1717296;
                12'd2068: exp <= 22'd1716296;
                12'd2069: exp <= 22'd1715295;
                12'd2070: exp <= 22'd1714295;
                12'd2071: exp <= 22'd1713296;
                12'd2072: exp <= 22'd1712296;
                12'd2073: exp <= 22'd1711297;
                12'd2074: exp <= 22'd1710297;
                12'd2075: exp <= 22'd1709298;
                12'd2076: exp <= 22'd1708299;
                12'd2077: exp <= 22'd1707300;
                12'd2078: exp <= 22'd1706302;
                12'd2079: exp <= 22'd1705303;
                12'd2080: exp <= 22'd1704305;
                12'd2081: exp <= 22'd1703307;
                12'd2082: exp <= 22'd1702309;
                12'd2083: exp <= 22'd1701311;
                12'd2084: exp <= 22'd1700314;
                12'd2085: exp <= 22'd1699316;
                12'd2086: exp <= 22'd1698319;
                12'd2087: exp <= 22'd1697322;
                12'd2088: exp <= 22'd1696325;
                12'd2089: exp <= 22'd1695328;
                12'd2090: exp <= 22'd1694332;
                12'd2091: exp <= 22'd1693335;
                12'd2092: exp <= 22'd1692339;
                12'd2093: exp <= 22'd1691343;
                12'd2094: exp <= 22'd1690347;
                12'd2095: exp <= 22'd1689351;
                12'd2096: exp <= 22'd1688356;
                12'd2097: exp <= 22'd1687360;
                12'd2098: exp <= 22'd1686365;
                12'd2099: exp <= 22'd1685370;
                12'd2100: exp <= 22'd1684375;
                12'd2101: exp <= 22'd1683380;
                12'd2102: exp <= 22'd1682386;
                12'd2103: exp <= 22'd1681391;
                12'd2104: exp <= 22'd1680397;
                12'd2105: exp <= 22'd1679403;
                12'd2106: exp <= 22'd1678409;
                12'd2107: exp <= 22'd1677415;
                12'd2108: exp <= 22'd1676422;
                12'd2109: exp <= 22'd1675428;
                12'd2110: exp <= 22'd1674435;
                12'd2111: exp <= 22'd1673442;
                12'd2112: exp <= 22'd1672449;
                12'd2113: exp <= 22'd1671456;
                12'd2114: exp <= 22'd1670464;
                12'd2115: exp <= 22'd1669471;
                12'd2116: exp <= 22'd1668479;
                12'd2117: exp <= 22'd1667487;
                12'd2118: exp <= 22'd1666495;
                12'd2119: exp <= 22'd1665504;
                12'd2120: exp <= 22'd1664512;
                12'd2121: exp <= 22'd1663521;
                12'd2122: exp <= 22'd1662530;
                12'd2123: exp <= 22'd1661538;
                12'd2124: exp <= 22'd1660548;
                12'd2125: exp <= 22'd1659557;
                12'd2126: exp <= 22'd1658566;
                12'd2127: exp <= 22'd1657576;
                12'd2128: exp <= 22'd1656586;
                12'd2129: exp <= 22'd1655596;
                12'd2130: exp <= 22'd1654606;
                12'd2131: exp <= 22'd1653616;
                12'd2132: exp <= 22'd1652627;
                12'd2133: exp <= 22'd1651637;
                12'd2134: exp <= 22'd1650648;
                12'd2135: exp <= 22'd1649659;
                12'd2136: exp <= 22'd1648670;
                12'd2137: exp <= 22'd1647681;
                12'd2138: exp <= 22'd1646693;
                12'd2139: exp <= 22'd1645705;
                12'd2140: exp <= 22'd1644716;
                12'd2141: exp <= 22'd1643728;
                12'd2142: exp <= 22'd1642741;
                12'd2143: exp <= 22'd1641753;
                12'd2144: exp <= 22'd1640765;
                12'd2145: exp <= 22'd1639778;
                12'd2146: exp <= 22'd1638791;
                12'd2147: exp <= 22'd1637804;
                12'd2148: exp <= 22'd1636817;
                12'd2149: exp <= 22'd1635830;
                12'd2150: exp <= 22'd1634844;
                12'd2151: exp <= 22'd1633857;
                12'd2152: exp <= 22'd1632871;
                12'd2153: exp <= 22'd1631885;
                12'd2154: exp <= 22'd1630899;
                12'd2155: exp <= 22'd1629914;
                12'd2156: exp <= 22'd1628928;
                12'd2157: exp <= 22'd1627943;
                12'd2158: exp <= 22'd1626957;
                12'd2159: exp <= 22'd1625972;
                12'd2160: exp <= 22'd1624988;
                12'd2161: exp <= 22'd1624003;
                12'd2162: exp <= 22'd1623018;
                12'd2163: exp <= 22'd1622034;
                12'd2164: exp <= 22'd1621050;
                12'd2165: exp <= 22'd1620066;
                12'd2166: exp <= 22'd1619082;
                12'd2167: exp <= 22'd1618098;
                12'd2168: exp <= 22'd1617115;
                12'd2169: exp <= 22'd1616131;
                12'd2170: exp <= 22'd1615148;
                12'd2171: exp <= 22'd1614165;
                12'd2172: exp <= 22'd1613182;
                12'd2173: exp <= 22'd1612200;
                12'd2174: exp <= 22'd1611217;
                12'd2175: exp <= 22'd1610235;
                12'd2176: exp <= 22'd1609253;
                12'd2177: exp <= 22'd1608271;
                12'd2178: exp <= 22'd1607289;
                12'd2179: exp <= 22'd1606307;
                12'd2180: exp <= 22'd1605325;
                12'd2181: exp <= 22'd1604344;
                12'd2182: exp <= 22'd1603363;
                12'd2183: exp <= 22'd1602382;
                12'd2184: exp <= 22'd1601401;
                12'd2185: exp <= 22'd1600420;
                12'd2186: exp <= 22'd1599440;
                12'd2187: exp <= 22'd1598459;
                12'd2188: exp <= 22'd1597479;
                12'd2189: exp <= 22'd1596499;
                12'd2190: exp <= 22'd1595519;
                12'd2191: exp <= 22'd1594540;
                12'd2192: exp <= 22'd1593560;
                12'd2193: exp <= 22'd1592581;
                12'd2194: exp <= 22'd1591601;
                12'd2195: exp <= 22'd1590622;
                12'd2196: exp <= 22'd1589644;
                12'd2197: exp <= 22'd1588665;
                12'd2198: exp <= 22'd1587686;
                12'd2199: exp <= 22'd1586708;
                12'd2200: exp <= 22'd1585730;
                12'd2201: exp <= 22'd1584752;
                12'd2202: exp <= 22'd1583774;
                12'd2203: exp <= 22'd1582796;
                12'd2204: exp <= 22'd1581819;
                12'd2205: exp <= 22'd1580841;
                12'd2206: exp <= 22'd1579864;
                12'd2207: exp <= 22'd1578887;
                12'd2208: exp <= 22'd1577910;
                12'd2209: exp <= 22'd1576933;
                12'd2210: exp <= 22'd1575957;
                12'd2211: exp <= 22'd1574980;
                12'd2212: exp <= 22'd1574004;
                12'd2213: exp <= 22'd1573028;
                12'd2214: exp <= 22'd1572052;
                12'd2215: exp <= 22'd1571076;
                12'd2216: exp <= 22'd1570101;
                12'd2217: exp <= 22'd1569125;
                12'd2218: exp <= 22'd1568150;
                12'd2219: exp <= 22'd1567175;
                12'd2220: exp <= 22'd1566200;
                12'd2221: exp <= 22'd1565226;
                12'd2222: exp <= 22'd1564251;
                12'd2223: exp <= 22'd1563277;
                12'd2224: exp <= 22'd1562302;
                12'd2225: exp <= 22'd1561328;
                12'd2226: exp <= 22'd1560354;
                12'd2227: exp <= 22'd1559381;
                12'd2228: exp <= 22'd1558407;
                12'd2229: exp <= 22'd1557434;
                12'd2230: exp <= 22'd1556460;
                12'd2231: exp <= 22'd1555487;
                12'd2232: exp <= 22'd1554514;
                12'd2233: exp <= 22'd1553541;
                12'd2234: exp <= 22'd1552569;
                12'd2235: exp <= 22'd1551596;
                12'd2236: exp <= 22'd1550624;
                12'd2237: exp <= 22'd1549652;
                12'd2238: exp <= 22'd1548680;
                12'd2239: exp <= 22'd1547708;
                12'd2240: exp <= 22'd1546737;
                12'd2241: exp <= 22'd1545765;
                12'd2242: exp <= 22'd1544794;
                12'd2243: exp <= 22'd1543823;
                12'd2244: exp <= 22'd1542852;
                12'd2245: exp <= 22'd1541881;
                12'd2246: exp <= 22'd1540911;
                12'd2247: exp <= 22'd1539940;
                12'd2248: exp <= 22'd1538970;
                12'd2249: exp <= 22'd1538000;
                12'd2250: exp <= 22'd1537030;
                12'd2251: exp <= 22'd1536060;
                12'd2252: exp <= 22'd1535090;
                12'd2253: exp <= 22'd1534121;
                12'd2254: exp <= 22'd1533151;
                12'd2255: exp <= 22'd1532182;
                12'd2256: exp <= 22'd1531213;
                12'd2257: exp <= 22'd1530244;
                12'd2258: exp <= 22'd1529276;
                12'd2259: exp <= 22'd1528307;
                12'd2260: exp <= 22'd1527339;
                12'd2261: exp <= 22'd1526371;
                12'd2262: exp <= 22'd1525403;
                12'd2263: exp <= 22'd1524435;
                12'd2264: exp <= 22'd1523467;
                12'd2265: exp <= 22'd1522500;
                12'd2266: exp <= 22'd1521532;
                12'd2267: exp <= 22'd1520565;
                12'd2268: exp <= 22'd1519598;
                12'd2269: exp <= 22'd1518631;
                12'd2270: exp <= 22'd1517665;
                12'd2271: exp <= 22'd1516698;
                12'd2272: exp <= 22'd1515732;
                12'd2273: exp <= 22'd1514766;
                12'd2274: exp <= 22'd1513800;
                12'd2275: exp <= 22'd1512834;
                12'd2276: exp <= 22'd1511868;
                12'd2277: exp <= 22'd1510902;
                12'd2278: exp <= 22'd1509937;
                12'd2279: exp <= 22'd1508972;
                12'd2280: exp <= 22'd1508007;
                12'd2281: exp <= 22'd1507042;
                12'd2282: exp <= 22'd1506077;
                12'd2283: exp <= 22'd1505113;
                12'd2284: exp <= 22'd1504148;
                12'd2285: exp <= 22'd1503184;
                12'd2286: exp <= 22'd1502220;
                12'd2287: exp <= 22'd1501256;
                12'd2288: exp <= 22'd1500292;
                12'd2289: exp <= 22'd1499329;
                12'd2290: exp <= 22'd1498365;
                12'd2291: exp <= 22'd1497402;
                12'd2292: exp <= 22'd1496439;
                12'd2293: exp <= 22'd1495476;
                12'd2294: exp <= 22'd1494513;
                12'd2295: exp <= 22'd1493550;
                12'd2296: exp <= 22'd1492588;
                12'd2297: exp <= 22'd1491626;
                12'd2298: exp <= 22'd1490664;
                12'd2299: exp <= 22'd1489702;
                12'd2300: exp <= 22'd1488740;
                12'd2301: exp <= 22'd1487778;
                12'd2302: exp <= 22'd1486817;
                12'd2303: exp <= 22'd1485855;
                12'd2304: exp <= 22'd1484894;
                12'd2305: exp <= 22'd1483933;
                12'd2306: exp <= 22'd1482973;
                12'd2307: exp <= 22'd1482012;
                12'd2308: exp <= 22'd1481051;
                12'd2309: exp <= 22'd1480091;
                12'd2310: exp <= 22'd1479131;
                12'd2311: exp <= 22'd1478171;
                12'd2312: exp <= 22'd1477211;
                12'd2313: exp <= 22'd1476251;
                12'd2314: exp <= 22'd1475292;
                12'd2315: exp <= 22'd1474332;
                12'd2316: exp <= 22'd1473373;
                12'd2317: exp <= 22'd1472414;
                12'd2318: exp <= 22'd1471455;
                12'd2319: exp <= 22'd1470497;
                12'd2320: exp <= 22'd1469538;
                12'd2321: exp <= 22'd1468580;
                12'd2322: exp <= 22'd1467621;
                12'd2323: exp <= 22'd1466663;
                12'd2324: exp <= 22'd1465706;
                12'd2325: exp <= 22'd1464748;
                12'd2326: exp <= 22'd1463790;
                12'd2327: exp <= 22'd1462833;
                12'd2328: exp <= 22'd1461876;
                12'd2329: exp <= 22'd1460918;
                12'd2330: exp <= 22'd1459962;
                12'd2331: exp <= 22'd1459005;
                12'd2332: exp <= 22'd1458048;
                12'd2333: exp <= 22'd1457092;
                12'd2334: exp <= 22'd1456135;
                12'd2335: exp <= 22'd1455179;
                12'd2336: exp <= 22'd1454223;
                12'd2337: exp <= 22'd1453268;
                12'd2338: exp <= 22'd1452312;
                12'd2339: exp <= 22'd1451356;
                12'd2340: exp <= 22'd1450401;
                12'd2341: exp <= 22'd1449446;
                12'd2342: exp <= 22'd1448491;
                12'd2343: exp <= 22'd1447536;
                12'd2344: exp <= 22'd1446582;
                12'd2345: exp <= 22'd1445627;
                12'd2346: exp <= 22'd1444673;
                12'd2347: exp <= 22'd1443719;
                12'd2348: exp <= 22'd1442765;
                12'd2349: exp <= 22'd1441811;
                12'd2350: exp <= 22'd1440857;
                12'd2351: exp <= 22'd1439903;
                12'd2352: exp <= 22'd1438950;
                12'd2353: exp <= 22'd1437997;
                12'd2354: exp <= 22'd1437044;
                12'd2355: exp <= 22'd1436091;
                12'd2356: exp <= 22'd1435138;
                12'd2357: exp <= 22'd1434186;
                12'd2358: exp <= 22'd1433233;
                12'd2359: exp <= 22'd1432281;
                12'd2360: exp <= 22'd1431329;
                12'd2361: exp <= 22'd1430377;
                12'd2362: exp <= 22'd1429425;
                12'd2363: exp <= 22'd1428474;
                12'd2364: exp <= 22'd1427522;
                12'd2365: exp <= 22'd1426571;
                12'd2366: exp <= 22'd1425620;
                12'd2367: exp <= 22'd1424669;
                12'd2368: exp <= 22'd1423718;
                12'd2369: exp <= 22'd1422767;
                12'd2370: exp <= 22'd1421817;
                12'd2371: exp <= 22'd1420867;
                12'd2372: exp <= 22'd1419917;
                12'd2373: exp <= 22'd1418967;
                12'd2374: exp <= 22'd1418017;
                12'd2375: exp <= 22'd1417067;
                12'd2376: exp <= 22'd1416118;
                12'd2377: exp <= 22'd1415168;
                12'd2378: exp <= 22'd1414219;
                12'd2379: exp <= 22'd1413270;
                12'd2380: exp <= 22'd1412321;
                12'd2381: exp <= 22'd1411372;
                12'd2382: exp <= 22'd1410424;
                12'd2383: exp <= 22'd1409475;
                12'd2384: exp <= 22'd1408527;
                12'd2385: exp <= 22'd1407579;
                12'd2386: exp <= 22'd1406631;
                12'd2387: exp <= 22'd1405684;
                12'd2388: exp <= 22'd1404736;
                12'd2389: exp <= 22'd1403789;
                12'd2390: exp <= 22'd1402841;
                12'd2391: exp <= 22'd1401894;
                12'd2392: exp <= 22'd1400947;
                12'd2393: exp <= 22'd1400000;
                12'd2394: exp <= 22'd1399054;
                12'd2395: exp <= 22'd1398107;
                12'd2396: exp <= 22'd1397161;
                12'd2397: exp <= 22'd1396215;
                12'd2398: exp <= 22'd1395269;
                12'd2399: exp <= 22'd1394323;
                12'd2400: exp <= 22'd1393378;
                12'd2401: exp <= 22'd1392432;
                12'd2402: exp <= 22'd1391487;
                12'd2403: exp <= 22'd1390541;
                12'd2404: exp <= 22'd1389596;
                12'd2405: exp <= 22'd1388652;
                12'd2406: exp <= 22'd1387707;
                12'd2407: exp <= 22'd1386762;
                12'd2408: exp <= 22'd1385818;
                12'd2409: exp <= 22'd1384874;
                12'd2410: exp <= 22'd1383930;
                12'd2411: exp <= 22'd1382986;
                12'd2412: exp <= 22'd1382042;
                12'd2413: exp <= 22'd1381099;
                12'd2414: exp <= 22'd1380155;
                12'd2415: exp <= 22'd1379212;
                12'd2416: exp <= 22'd1378269;
                12'd2417: exp <= 22'd1377326;
                12'd2418: exp <= 22'd1376383;
                12'd2419: exp <= 22'd1375440;
                12'd2420: exp <= 22'd1374498;
                12'd2421: exp <= 22'd1373556;
                12'd2422: exp <= 22'd1372613;
                12'd2423: exp <= 22'd1371671;
                12'd2424: exp <= 22'd1370730;
                12'd2425: exp <= 22'd1369788;
                12'd2426: exp <= 22'd1368846;
                12'd2427: exp <= 22'd1367905;
                12'd2428: exp <= 22'd1366964;
                12'd2429: exp <= 22'd1366023;
                12'd2430: exp <= 22'd1365082;
                12'd2431: exp <= 22'd1364141;
                12'd2432: exp <= 22'd1363201;
                12'd2433: exp <= 22'd1362260;
                12'd2434: exp <= 22'd1361320;
                12'd2435: exp <= 22'd1360380;
                12'd2436: exp <= 22'd1359440;
                12'd2437: exp <= 22'd1358500;
                12'd2438: exp <= 22'd1357561;
                12'd2439: exp <= 22'd1356621;
                12'd2440: exp <= 22'd1355682;
                12'd2441: exp <= 22'd1354743;
                12'd2442: exp <= 22'd1353804;
                12'd2443: exp <= 22'd1352865;
                12'd2444: exp <= 22'd1351927;
                12'd2445: exp <= 22'd1350988;
                12'd2446: exp <= 22'd1350050;
                12'd2447: exp <= 22'd1349112;
                12'd2448: exp <= 22'd1348174;
                12'd2449: exp <= 22'd1347236;
                12'd2450: exp <= 22'd1346298;
                12'd2451: exp <= 22'd1345361;
                12'd2452: exp <= 22'd1344423;
                12'd2453: exp <= 22'd1343486;
                12'd2454: exp <= 22'd1342549;
                12'd2455: exp <= 22'd1341612;
                12'd2456: exp <= 22'd1340675;
                12'd2457: exp <= 22'd1339739;
                12'd2458: exp <= 22'd1338802;
                12'd2459: exp <= 22'd1337866;
                12'd2460: exp <= 22'd1336930;
                12'd2461: exp <= 22'd1335994;
                12'd2462: exp <= 22'd1335058;
                12'd2463: exp <= 22'd1334123;
                12'd2464: exp <= 22'd1333187;
                12'd2465: exp <= 22'd1332252;
                12'd2466: exp <= 22'd1331317;
                12'd2467: exp <= 22'd1330382;
                12'd2468: exp <= 22'd1329447;
                12'd2469: exp <= 22'd1328512;
                12'd2470: exp <= 22'd1327578;
                12'd2471: exp <= 22'd1326643;
                12'd2472: exp <= 22'd1325709;
                12'd2473: exp <= 22'd1324775;
                12'd2474: exp <= 22'd1323841;
                12'd2475: exp <= 22'd1322907;
                12'd2476: exp <= 22'd1321974;
                12'd2477: exp <= 22'd1321040;
                12'd2478: exp <= 22'd1320107;
                12'd2479: exp <= 22'd1319174;
                12'd2480: exp <= 22'd1318241;
                12'd2481: exp <= 22'd1317308;
                12'd2482: exp <= 22'd1316376;
                12'd2483: exp <= 22'd1315443;
                12'd2484: exp <= 22'd1314511;
                12'd2485: exp <= 22'd1313579;
                12'd2486: exp <= 22'd1312647;
                12'd2487: exp <= 22'd1311715;
                12'd2488: exp <= 22'd1310783;
                12'd2489: exp <= 22'd1309852;
                12'd2490: exp <= 22'd1308920;
                12'd2491: exp <= 22'd1307989;
                12'd2492: exp <= 22'd1307058;
                12'd2493: exp <= 22'd1306127;
                12'd2494: exp <= 22'd1305196;
                12'd2495: exp <= 22'd1304266;
                12'd2496: exp <= 22'd1303335;
                12'd2497: exp <= 22'd1302405;
                12'd2498: exp <= 22'd1301475;
                12'd2499: exp <= 22'd1300545;
                12'd2500: exp <= 22'd1299615;
                12'd2501: exp <= 22'd1298686;
                12'd2502: exp <= 22'd1297756;
                12'd2503: exp <= 22'd1296827;
                12'd2504: exp <= 22'd1295898;
                12'd2505: exp <= 22'd1294969;
                12'd2506: exp <= 22'd1294040;
                12'd2507: exp <= 22'd1293111;
                12'd2508: exp <= 22'd1292183;
                12'd2509: exp <= 22'd1291254;
                12'd2510: exp <= 22'd1290326;
                12'd2511: exp <= 22'd1289398;
                12'd2512: exp <= 22'd1288470;
                12'd2513: exp <= 22'd1287542;
                12'd2514: exp <= 22'd1286615;
                12'd2515: exp <= 22'd1285687;
                12'd2516: exp <= 22'd1284760;
                12'd2517: exp <= 22'd1283833;
                12'd2518: exp <= 22'd1282906;
                12'd2519: exp <= 22'd1281979;
                12'd2520: exp <= 22'd1281053;
                12'd2521: exp <= 22'd1280126;
                12'd2522: exp <= 22'd1279200;
                12'd2523: exp <= 22'd1278274;
                12'd2524: exp <= 22'd1277348;
                12'd2525: exp <= 22'd1276422;
                12'd2526: exp <= 22'd1275496;
                12'd2527: exp <= 22'd1274570;
                12'd2528: exp <= 22'd1273645;
                12'd2529: exp <= 22'd1272720;
                12'd2530: exp <= 22'd1271795;
                12'd2531: exp <= 22'd1270870;
                12'd2532: exp <= 22'd1269945;
                12'd2533: exp <= 22'd1269020;
                12'd2534: exp <= 22'd1268096;
                12'd2535: exp <= 22'd1267172;
                12'd2536: exp <= 22'd1266247;
                12'd2537: exp <= 22'd1265324;
                12'd2538: exp <= 22'd1264400;
                12'd2539: exp <= 22'd1263476;
                12'd2540: exp <= 22'd1262552;
                12'd2541: exp <= 22'd1261629;
                12'd2542: exp <= 22'd1260706;
                12'd2543: exp <= 22'd1259783;
                12'd2544: exp <= 22'd1258860;
                12'd2545: exp <= 22'd1257937;
                12'd2546: exp <= 22'd1257015;
                12'd2547: exp <= 22'd1256092;
                12'd2548: exp <= 22'd1255170;
                12'd2549: exp <= 22'd1254248;
                12'd2550: exp <= 22'd1253326;
                12'd2551: exp <= 22'd1252404;
                12'd2552: exp <= 22'd1251482;
                12'd2553: exp <= 22'd1250561;
                12'd2554: exp <= 22'd1249640;
                12'd2555: exp <= 22'd1248718;
                12'd2556: exp <= 22'd1247797;
                12'd2557: exp <= 22'd1246877;
                12'd2558: exp <= 22'd1245956;
                12'd2559: exp <= 22'd1245035;
                12'd2560: exp <= 22'd1244115;
                12'd2561: exp <= 22'd1243195;
                12'd2562: exp <= 22'd1242275;
                12'd2563: exp <= 22'd1241355;
                12'd2564: exp <= 22'd1240435;
                12'd2565: exp <= 22'd1239515;
                12'd2566: exp <= 22'd1238596;
                12'd2567: exp <= 22'd1237677;
                12'd2568: exp <= 22'd1236757;
                12'd2569: exp <= 22'd1235838;
                12'd2570: exp <= 22'd1234920;
                12'd2571: exp <= 22'd1234001;
                12'd2572: exp <= 22'd1233082;
                12'd2573: exp <= 22'd1232164;
                12'd2574: exp <= 22'd1231246;
                12'd2575: exp <= 22'd1230328;
                12'd2576: exp <= 22'd1229410;
                12'd2577: exp <= 22'd1228492;
                12'd2578: exp <= 22'd1227574;
                12'd2579: exp <= 22'd1226657;
                12'd2580: exp <= 22'd1225740;
                12'd2581: exp <= 22'd1224823;
                12'd2582: exp <= 22'd1223906;
                12'd2583: exp <= 22'd1222989;
                12'd2584: exp <= 22'd1222072;
                12'd2585: exp <= 22'd1221156;
                12'd2586: exp <= 22'd1220239;
                12'd2587: exp <= 22'd1219323;
                12'd2588: exp <= 22'd1218407;
                12'd2589: exp <= 22'd1217491;
                12'd2590: exp <= 22'd1216575;
                12'd2591: exp <= 22'd1215660;
                12'd2592: exp <= 22'd1214744;
                12'd2593: exp <= 22'd1213829;
                12'd2594: exp <= 22'd1212914;
                12'd2595: exp <= 22'd1211999;
                12'd2596: exp <= 22'd1211084;
                12'd2597: exp <= 22'd1210170;
                12'd2598: exp <= 22'd1209255;
                12'd2599: exp <= 22'd1208341;
                12'd2600: exp <= 22'd1207427;
                12'd2601: exp <= 22'd1206512;
                12'd2602: exp <= 22'd1205599;
                12'd2603: exp <= 22'd1204685;
                12'd2604: exp <= 22'd1203771;
                12'd2605: exp <= 22'd1202858;
                12'd2606: exp <= 22'd1201945;
                12'd2607: exp <= 22'd1201032;
                12'd2608: exp <= 22'd1200119;
                12'd2609: exp <= 22'd1199206;
                12'd2610: exp <= 22'd1198293;
                12'd2611: exp <= 22'd1197381;
                12'd2612: exp <= 22'd1196468;
                12'd2613: exp <= 22'd1195556;
                12'd2614: exp <= 22'd1194644;
                12'd2615: exp <= 22'd1193732;
                12'd2616: exp <= 22'd1192821;
                12'd2617: exp <= 22'd1191909;
                12'd2618: exp <= 22'd1190998;
                12'd2619: exp <= 22'd1190086;
                12'd2620: exp <= 22'd1189175;
                12'd2621: exp <= 22'd1188264;
                12'd2622: exp <= 22'd1187353;
                12'd2623: exp <= 22'd1186443;
                12'd2624: exp <= 22'd1185532;
                12'd2625: exp <= 22'd1184622;
                12'd2626: exp <= 22'd1183712;
                12'd2627: exp <= 22'd1182802;
                12'd2628: exp <= 22'd1181892;
                12'd2629: exp <= 22'd1180982;
                12'd2630: exp <= 22'd1180073;
                12'd2631: exp <= 22'd1179163;
                12'd2632: exp <= 22'd1178254;
                12'd2633: exp <= 22'd1177345;
                12'd2634: exp <= 22'd1176436;
                12'd2635: exp <= 22'd1175527;
                12'd2636: exp <= 22'd1174619;
                12'd2637: exp <= 22'd1173710;
                12'd2638: exp <= 22'd1172802;
                12'd2639: exp <= 22'd1171894;
                12'd2640: exp <= 22'd1170986;
                12'd2641: exp <= 22'd1170078;
                12'd2642: exp <= 22'd1169170;
                12'd2643: exp <= 22'd1168262;
                12'd2644: exp <= 22'd1167355;
                12'd2645: exp <= 22'd1166448;
                12'd2646: exp <= 22'd1165541;
                12'd2647: exp <= 22'd1164634;
                12'd2648: exp <= 22'd1163727;
                12'd2649: exp <= 22'd1162820;
                12'd2650: exp <= 22'd1161914;
                12'd2651: exp <= 22'd1161007;
                12'd2652: exp <= 22'd1160101;
                12'd2653: exp <= 22'd1159195;
                12'd2654: exp <= 22'd1158289;
                12'd2655: exp <= 22'd1157384;
                12'd2656: exp <= 22'd1156478;
                12'd2657: exp <= 22'd1155573;
                12'd2658: exp <= 22'd1154667;
                12'd2659: exp <= 22'd1153762;
                12'd2660: exp <= 22'd1152857;
                12'd2661: exp <= 22'd1151953;
                12'd2662: exp <= 22'd1151048;
                12'd2663: exp <= 22'd1150143;
                12'd2664: exp <= 22'd1149239;
                12'd2665: exp <= 22'd1148335;
                12'd2666: exp <= 22'd1147431;
                12'd2667: exp <= 22'd1146527;
                12'd2668: exp <= 22'd1145623;
                12'd2669: exp <= 22'd1144720;
                12'd2670: exp <= 22'd1143816;
                12'd2671: exp <= 22'd1142913;
                12'd2672: exp <= 22'd1142010;
                12'd2673: exp <= 22'd1141107;
                12'd2674: exp <= 22'd1140204;
                12'd2675: exp <= 22'd1139301;
                12'd2676: exp <= 22'd1138399;
                12'd2677: exp <= 22'd1137497;
                12'd2678: exp <= 22'd1136594;
                12'd2679: exp <= 22'd1135692;
                12'd2680: exp <= 22'd1134790;
                12'd2681: exp <= 22'd1133889;
                12'd2682: exp <= 22'd1132987;
                12'd2683: exp <= 22'd1132086;
                12'd2684: exp <= 22'd1131184;
                12'd2685: exp <= 22'd1130283;
                12'd2686: exp <= 22'd1129382;
                12'd2687: exp <= 22'd1128482;
                12'd2688: exp <= 22'd1127581;
                12'd2689: exp <= 22'd1126680;
                12'd2690: exp <= 22'd1125780;
                12'd2691: exp <= 22'd1124880;
                12'd2692: exp <= 22'd1123980;
                12'd2693: exp <= 22'd1123080;
                12'd2694: exp <= 22'd1122180;
                12'd2695: exp <= 22'd1121280;
                12'd2696: exp <= 22'd1120381;
                12'd2697: exp <= 22'd1119482;
                12'd2698: exp <= 22'd1118582;
                12'd2699: exp <= 22'd1117683;
                12'd2700: exp <= 22'd1116785;
                12'd2701: exp <= 22'd1115886;
                12'd2702: exp <= 22'd1114987;
                12'd2703: exp <= 22'd1114089;
                12'd2704: exp <= 22'd1113191;
                12'd2705: exp <= 22'd1112293;
                12'd2706: exp <= 22'd1111395;
                12'd2707: exp <= 22'd1110497;
                12'd2708: exp <= 22'd1109599;
                12'd2709: exp <= 22'd1108702;
                12'd2710: exp <= 22'd1107805;
                12'd2711: exp <= 22'd1106907;
                12'd2712: exp <= 22'd1106010;
                12'd2713: exp <= 22'd1105113;
                12'd2714: exp <= 22'd1104217;
                12'd2715: exp <= 22'd1103320;
                12'd2716: exp <= 22'd1102424;
                12'd2717: exp <= 22'd1101527;
                12'd2718: exp <= 22'd1100631;
                12'd2719: exp <= 22'd1099735;
                12'd2720: exp <= 22'd1098840;
                12'd2721: exp <= 22'd1097944;
                12'd2722: exp <= 22'd1097048;
                12'd2723: exp <= 22'd1096153;
                12'd2724: exp <= 22'd1095258;
                12'd2725: exp <= 22'd1094363;
                12'd2726: exp <= 22'd1093468;
                12'd2727: exp <= 22'd1092573;
                12'd2728: exp <= 22'd1091679;
                12'd2729: exp <= 22'd1090784;
                12'd2730: exp <= 22'd1089890;
                12'd2731: exp <= 22'd1088996;
                12'd2732: exp <= 22'd1088102;
                12'd2733: exp <= 22'd1087208;
                12'd2734: exp <= 22'd1086314;
                12'd2735: exp <= 22'd1085421;
                12'd2736: exp <= 22'd1084527;
                12'd2737: exp <= 22'd1083634;
                12'd2738: exp <= 22'd1082741;
                12'd2739: exp <= 22'd1081848;
                12'd2740: exp <= 22'd1080955;
                12'd2741: exp <= 22'd1080063;
                12'd2742: exp <= 22'd1079170;
                12'd2743: exp <= 22'd1078278;
                12'd2744: exp <= 22'd1077386;
                12'd2745: exp <= 22'd1076494;
                12'd2746: exp <= 22'd1075602;
                12'd2747: exp <= 22'd1074710;
                12'd2748: exp <= 22'd1073818;
                12'd2749: exp <= 22'd1072927;
                12'd2750: exp <= 22'd1072036;
                12'd2751: exp <= 22'd1071145;
                12'd2752: exp <= 22'd1070254;
                12'd2753: exp <= 22'd1069363;
                12'd2754: exp <= 22'd1068472;
                12'd2755: exp <= 22'd1067582;
                12'd2756: exp <= 22'd1066691;
                12'd2757: exp <= 22'd1065801;
                12'd2758: exp <= 22'd1064911;
                12'd2759: exp <= 22'd1064021;
                12'd2760: exp <= 22'd1063131;
                12'd2761: exp <= 22'd1062242;
                12'd2762: exp <= 22'd1061352;
                12'd2763: exp <= 22'd1060463;
                12'd2764: exp <= 22'd1059574;
                12'd2765: exp <= 22'd1058685;
                12'd2766: exp <= 22'd1057796;
                12'd2767: exp <= 22'd1056907;
                12'd2768: exp <= 22'd1056018;
                12'd2769: exp <= 22'd1055130;
                12'd2770: exp <= 22'd1054242;
                12'd2771: exp <= 22'd1053354;
                12'd2772: exp <= 22'd1052466;
                12'd2773: exp <= 22'd1051578;
                12'd2774: exp <= 22'd1050690;
                12'd2775: exp <= 22'd1049803;
                12'd2776: exp <= 22'd1048915;
                12'd2777: exp <= 22'd1048028;
                12'd2778: exp <= 22'd1047141;
                12'd2779: exp <= 22'd1046254;
                12'd2780: exp <= 22'd1045367;
                12'd2781: exp <= 22'd1044481;
                12'd2782: exp <= 22'd1043594;
                12'd2783: exp <= 22'd1042708;
                12'd2784: exp <= 22'd1041822;
                12'd2785: exp <= 22'd1040936;
                12'd2786: exp <= 22'd1040050;
                12'd2787: exp <= 22'd1039164;
                12'd2788: exp <= 22'd1038279;
                12'd2789: exp <= 22'd1037393;
                12'd2790: exp <= 22'd1036508;
                12'd2791: exp <= 22'd1035623;
                12'd2792: exp <= 22'd1034738;
                12'd2793: exp <= 22'd1033853;
                12'd2794: exp <= 22'd1032969;
                12'd2795: exp <= 22'd1032084;
                12'd2796: exp <= 22'd1031200;
                12'd2797: exp <= 22'd1030315;
                12'd2798: exp <= 22'd1029431;
                12'd2799: exp <= 22'd1028547;
                12'd2800: exp <= 22'd1027664;
                12'd2801: exp <= 22'd1026780;
                12'd2802: exp <= 22'd1025897;
                12'd2803: exp <= 22'd1025013;
                12'd2804: exp <= 22'd1024130;
                12'd2805: exp <= 22'd1023247;
                12'd2806: exp <= 22'd1022364;
                12'd2807: exp <= 22'd1021482;
                12'd2808: exp <= 22'd1020599;
                12'd2809: exp <= 22'd1019717;
                12'd2810: exp <= 22'd1018834;
                12'd2811: exp <= 22'd1017952;
                12'd2812: exp <= 22'd1017070;
                12'd2813: exp <= 22'd1016188;
                12'd2814: exp <= 22'd1015307;
                12'd2815: exp <= 22'd1014425;
                12'd2816: exp <= 22'd1013544;
                12'd2817: exp <= 22'd1012663;
                12'd2818: exp <= 22'd1011782;
                12'd2819: exp <= 22'd1010901;
                12'd2820: exp <= 22'd1010020;
                12'd2821: exp <= 22'd1009139;
                12'd2822: exp <= 22'd1008259;
                12'd2823: exp <= 22'd1007378;
                12'd2824: exp <= 22'd1006498;
                12'd2825: exp <= 22'd1005618;
                12'd2826: exp <= 22'd1004738;
                12'd2827: exp <= 22'd1003859;
                12'd2828: exp <= 22'd1002979;
                12'd2829: exp <= 22'd1002100;
                12'd2830: exp <= 22'd1001220;
                12'd2831: exp <= 22'd1000341;
                12'd2832: exp <= 22'd0999462;
                12'd2833: exp <= 22'd0998583;
                12'd2834: exp <= 22'd0997705;
                12'd2835: exp <= 22'd0996826;
                12'd2836: exp <= 22'd0995948;
                12'd2837: exp <= 22'd0995069;
                12'd2838: exp <= 22'd0994191;
                12'd2839: exp <= 22'd0993313;
                12'd2840: exp <= 22'd0992436;
                12'd2841: exp <= 22'd0991558;
                12'd2842: exp <= 22'd0990680;
                12'd2843: exp <= 22'd0989803;
                12'd2844: exp <= 22'd0988926;
                12'd2845: exp <= 22'd0988049;
                12'd2846: exp <= 22'd0987172;
                12'd2847: exp <= 22'd0986295;
                12'd2848: exp <= 22'd0985418;
                12'd2849: exp <= 22'd0984542;
                12'd2850: exp <= 22'd0983666;
                12'd2851: exp <= 22'd0982789;
                12'd2852: exp <= 22'd0981913;
                12'd2853: exp <= 22'd0981038;
                12'd2854: exp <= 22'd0980162;
                12'd2855: exp <= 22'd0979286;
                12'd2856: exp <= 22'd0978411;
                12'd2857: exp <= 22'd0977536;
                12'd2858: exp <= 22'd0976660;
                12'd2859: exp <= 22'd0975785;
                12'd2860: exp <= 22'd0974911;
                12'd2861: exp <= 22'd0974036;
                12'd2862: exp <= 22'd0973161;
                12'd2863: exp <= 22'd0972287;
                12'd2864: exp <= 22'd0971413;
                12'd2865: exp <= 22'd0970539;
                12'd2866: exp <= 22'd0969665;
                12'd2867: exp <= 22'd0968791;
                12'd2868: exp <= 22'd0967917;
                12'd2869: exp <= 22'd0967044;
                12'd2870: exp <= 22'd0966170;
                12'd2871: exp <= 22'd0965297;
                12'd2872: exp <= 22'd0964424;
                12'd2873: exp <= 22'd0963551;
                12'd2874: exp <= 22'd0962678;
                12'd2875: exp <= 22'd0961806;
                12'd2876: exp <= 22'd0960933;
                12'd2877: exp <= 22'd0960061;
                12'd2878: exp <= 22'd0959189;
                12'd2879: exp <= 22'd0958317;
                12'd2880: exp <= 22'd0957445;
                12'd2881: exp <= 22'd0956573;
                12'd2882: exp <= 22'd0955702;
                12'd2883: exp <= 22'd0954830;
                12'd2884: exp <= 22'd0953959;
                12'd2885: exp <= 22'd0953088;
                12'd2886: exp <= 22'd0952217;
                12'd2887: exp <= 22'd0951346;
                12'd2888: exp <= 22'd0950475;
                12'd2889: exp <= 22'd0949605;
                12'd2890: exp <= 22'd0948734;
                12'd2891: exp <= 22'd0947864;
                12'd2892: exp <= 22'd0946994;
                12'd2893: exp <= 22'd0946124;
                12'd2894: exp <= 22'd0945254;
                12'd2895: exp <= 22'd0944384;
                12'd2896: exp <= 22'd0943515;
                12'd2897: exp <= 22'd0942646;
                12'd2898: exp <= 22'd0941776;
                12'd2899: exp <= 22'd0940907;
                12'd2900: exp <= 22'd0940038;
                12'd2901: exp <= 22'd0939169;
                12'd2902: exp <= 22'd0938301;
                12'd2903: exp <= 22'd0937432;
                12'd2904: exp <= 22'd0936564;
                12'd2905: exp <= 22'd0935696;
                12'd2906: exp <= 22'd0934828;
                12'd2907: exp <= 22'd0933960;
                12'd2908: exp <= 22'd0933092;
                12'd2909: exp <= 22'd0932224;
                12'd2910: exp <= 22'd0931357;
                12'd2911: exp <= 22'd0930490;
                12'd2912: exp <= 22'd0929623;
                12'd2913: exp <= 22'd0928756;
                12'd2914: exp <= 22'd0927889;
                12'd2915: exp <= 22'd0927022;
                12'd2916: exp <= 22'd0926155;
                12'd2917: exp <= 22'd0925289;
                12'd2918: exp <= 22'd0924423;
                12'd2919: exp <= 22'd0923556;
                12'd2920: exp <= 22'd0922690;
                12'd2921: exp <= 22'd0921825;
                12'd2922: exp <= 22'd0920959;
                12'd2923: exp <= 22'd0920093;
                12'd2924: exp <= 22'd0919228;
                12'd2925: exp <= 22'd0918363;
                12'd2926: exp <= 22'd0917498;
                12'd2927: exp <= 22'd0916633;
                12'd2928: exp <= 22'd0915768;
                12'd2929: exp <= 22'd0914903;
                12'd2930: exp <= 22'd0914039;
                12'd2931: exp <= 22'd0913174;
                12'd2932: exp <= 22'd0912310;
                12'd2933: exp <= 22'd0911446;
                12'd2934: exp <= 22'd0910582;
                12'd2935: exp <= 22'd0909718;
                12'd2936: exp <= 22'd0908854;
                12'd2937: exp <= 22'd0907991;
                12'd2938: exp <= 22'd0907127;
                12'd2939: exp <= 22'd0906264;
                12'd2940: exp <= 22'd0905401;
                12'd2941: exp <= 22'd0904538;
                12'd2942: exp <= 22'd0903675;
                12'd2943: exp <= 22'd0902813;
                12'd2944: exp <= 22'd0901950;
                12'd2945: exp <= 22'd0901088;
                12'd2946: exp <= 22'd0900226;
                12'd2947: exp <= 22'd0899364;
                12'd2948: exp <= 22'd0898502;
                12'd2949: exp <= 22'd0897640;
                12'd2950: exp <= 22'd0896779;
                12'd2951: exp <= 22'd0895917;
                12'd2952: exp <= 22'd0895056;
                12'd2953: exp <= 22'd0894195;
                12'd2954: exp <= 22'd0893334;
                12'd2955: exp <= 22'd0892473;
                12'd2956: exp <= 22'd0891612;
                12'd2957: exp <= 22'd0890751;
                12'd2958: exp <= 22'd0889891;
                12'd2959: exp <= 22'd0889031;
                12'd2960: exp <= 22'd0888170;
                12'd2961: exp <= 22'd0887310;
                12'd2962: exp <= 22'd0886451;
                12'd2963: exp <= 22'd0885591;
                12'd2964: exp <= 22'd0884731;
                12'd2965: exp <= 22'd0883872;
                12'd2966: exp <= 22'd0883013;
                12'd2967: exp <= 22'd0882153;
                12'd2968: exp <= 22'd0881294;
                12'd2969: exp <= 22'd0880436;
                12'd2970: exp <= 22'd0879577;
                12'd2971: exp <= 22'd0878718;
                12'd2972: exp <= 22'd0877860;
                12'd2973: exp <= 22'd0877002;
                12'd2974: exp <= 22'd0876143;
                12'd2975: exp <= 22'd0875285;
                12'd2976: exp <= 22'd0874428;
                12'd2977: exp <= 22'd0873570;
                12'd2978: exp <= 22'd0872712;
                12'd2979: exp <= 22'd0871855;
                12'd2980: exp <= 22'd0870998;
                12'd2981: exp <= 22'd0870141;
                12'd2982: exp <= 22'd0869284;
                12'd2983: exp <= 22'd0868427;
                12'd2984: exp <= 22'd0867570;
                12'd2985: exp <= 22'd0866714;
                12'd2986: exp <= 22'd0865857;
                12'd2987: exp <= 22'd0865001;
                12'd2988: exp <= 22'd0864145;
                12'd2989: exp <= 22'd0863289;
                12'd2990: exp <= 22'd0862433;
                12'd2991: exp <= 22'd0861578;
                12'd2992: exp <= 22'd0860722;
                12'd2993: exp <= 22'd0859867;
                12'd2994: exp <= 22'd0859012;
                12'd2995: exp <= 22'd0858156;
                12'd2996: exp <= 22'd0857301;
                12'd2997: exp <= 22'd0856447;
                12'd2998: exp <= 22'd0855592;
                12'd2999: exp <= 22'd0854738;
                12'd3000: exp <= 22'd0853883;
                12'd3001: exp <= 22'd0853029;
                12'd3002: exp <= 22'd0852175;
                12'd3003: exp <= 22'd0851321;
                12'd3004: exp <= 22'd0850467;
                12'd3005: exp <= 22'd0849614;
                12'd3006: exp <= 22'd0848760;
                12'd3007: exp <= 22'd0847907;
                12'd3008: exp <= 22'd0847054;
                12'd3009: exp <= 22'd0846201;
                12'd3010: exp <= 22'd0845348;
                12'd3011: exp <= 22'd0844495;
                12'd3012: exp <= 22'd0843642;
                12'd3013: exp <= 22'd0842790;
                12'd3014: exp <= 22'd0841937;
                12'd3015: exp <= 22'd0841085;
                12'd3016: exp <= 22'd0840233;
                12'd3017: exp <= 22'd0839381;
                12'd3018: exp <= 22'd0838530;
                12'd3019: exp <= 22'd0837678;
                12'd3020: exp <= 22'd0836826;
                12'd3021: exp <= 22'd0835975;
                12'd3022: exp <= 22'd0835124;
                12'd3023: exp <= 22'd0834273;
                12'd3024: exp <= 22'd0833422;
                12'd3025: exp <= 22'd0832571;
                12'd3026: exp <= 22'd0831721;
                12'd3027: exp <= 22'd0830870;
                12'd3028: exp <= 22'd0830020;
                12'd3029: exp <= 22'd0829170;
                12'd3030: exp <= 22'd0828320;
                12'd3031: exp <= 22'd0827470;
                12'd3032: exp <= 22'd0826620;
                12'd3033: exp <= 22'd0825770;
                12'd3034: exp <= 22'd0824921;
                12'd3035: exp <= 22'd0824072;
                12'd3036: exp <= 22'd0823223;
                12'd3037: exp <= 22'd0822374;
                12'd3038: exp <= 22'd0821525;
                12'd3039: exp <= 22'd0820676;
                12'd3040: exp <= 22'd0819827;
                12'd3041: exp <= 22'd0818979;
                12'd3042: exp <= 22'd0818131;
                12'd3043: exp <= 22'd0817282;
                12'd3044: exp <= 22'd0816434;
                12'd3045: exp <= 22'd0815587;
                12'd3046: exp <= 22'd0814739;
                12'd3047: exp <= 22'd0813891;
                12'd3048: exp <= 22'd0813044;
                12'd3049: exp <= 22'd0812196;
                12'd3050: exp <= 22'd0811349;
                12'd3051: exp <= 22'd0810502;
                12'd3052: exp <= 22'd0809655;
                12'd3053: exp <= 22'd0808809;
                12'd3054: exp <= 22'd0807962;
                12'd3055: exp <= 22'd0807116;
                12'd3056: exp <= 22'd0806269;
                12'd3057: exp <= 22'd0805423;
                12'd3058: exp <= 22'd0804577;
                12'd3059: exp <= 22'd0803731;
                12'd3060: exp <= 22'd0802886;
                12'd3061: exp <= 22'd0802040;
                12'd3062: exp <= 22'd0801195;
                12'd3063: exp <= 22'd0800349;
                12'd3064: exp <= 22'd0799504;
                12'd3065: exp <= 22'd0798659;
                12'd3066: exp <= 22'd0797814;
                12'd3067: exp <= 22'd0796970;
                12'd3068: exp <= 22'd0796125;
                12'd3069: exp <= 22'd0795281;
                12'd3070: exp <= 22'd0794436;
                12'd3071: exp <= 22'd0793592;
                12'd3072: exp <= 22'd0792748;
                12'd3073: exp <= 22'd0791904;
                12'd3074: exp <= 22'd0791061;
                12'd3075: exp <= 22'd0790217;
                12'd3076: exp <= 22'd0789374;
                12'd3077: exp <= 22'd0788530;
                12'd3078: exp <= 22'd0787687;
                12'd3079: exp <= 22'd0786844;
                12'd3080: exp <= 22'd0786001;
                12'd3081: exp <= 22'd0785159;
                12'd3082: exp <= 22'd0784316;
                12'd3083: exp <= 22'd0783473;
                12'd3084: exp <= 22'd0782631;
                12'd3085: exp <= 22'd0781789;
                12'd3086: exp <= 22'd0780947;
                12'd3087: exp <= 22'd0780105;
                12'd3088: exp <= 22'd0779263;
                12'd3089: exp <= 22'd0778422;
                12'd3090: exp <= 22'd0777580;
                12'd3091: exp <= 22'd0776739;
                12'd3092: exp <= 22'd0775898;
                12'd3093: exp <= 22'd0775057;
                12'd3094: exp <= 22'd0774216;
                12'd3095: exp <= 22'd0773375;
                12'd3096: exp <= 22'd0772535;
                12'd3097: exp <= 22'd0771694;
                12'd3098: exp <= 22'd0770854;
                12'd3099: exp <= 22'd0770014;
                12'd3100: exp <= 22'd0769174;
                12'd3101: exp <= 22'd0768334;
                12'd3102: exp <= 22'd0767494;
                12'd3103: exp <= 22'd0766655;
                12'd3104: exp <= 22'd0765815;
                12'd3105: exp <= 22'd0764976;
                12'd3106: exp <= 22'd0764137;
                12'd3107: exp <= 22'd0763298;
                12'd3108: exp <= 22'd0762459;
                12'd3109: exp <= 22'd0761620;
                12'd3110: exp <= 22'd0760781;
                12'd3111: exp <= 22'd0759943;
                12'd3112: exp <= 22'd0759105;
                12'd3113: exp <= 22'd0758267;
                12'd3114: exp <= 22'd0757429;
                12'd3115: exp <= 22'd0756591;
                12'd3116: exp <= 22'd0755753;
                12'd3117: exp <= 22'd0754915;
                12'd3118: exp <= 22'd0754078;
                12'd3119: exp <= 22'd0753240;
                12'd3120: exp <= 22'd0752403;
                12'd3121: exp <= 22'd0751566;
                12'd3122: exp <= 22'd0750729;
                12'd3123: exp <= 22'd0749893;
                12'd3124: exp <= 22'd0749056;
                12'd3125: exp <= 22'd0748220;
                12'd3126: exp <= 22'd0747383;
                12'd3127: exp <= 22'd0746547;
                12'd3128: exp <= 22'd0745711;
                12'd3129: exp <= 22'd0744875;
                12'd3130: exp <= 22'd0744039;
                12'd3131: exp <= 22'd0743204;
                12'd3132: exp <= 22'd0742368;
                12'd3133: exp <= 22'd0741533;
                12'd3134: exp <= 22'd0740698;
                12'd3135: exp <= 22'd0739863;
                12'd3136: exp <= 22'd0739028;
                12'd3137: exp <= 22'd0738193;
                12'd3138: exp <= 22'd0737358;
                12'd3139: exp <= 22'd0736524;
                12'd3140: exp <= 22'd0735689;
                12'd3141: exp <= 22'd0734855;
                12'd3142: exp <= 22'd0734021;
                12'd3143: exp <= 22'd0733187;
                12'd3144: exp <= 22'd0732353;
                12'd3145: exp <= 22'd0731520;
                12'd3146: exp <= 22'd0730686;
                12'd3147: exp <= 22'd0729853;
                12'd3148: exp <= 22'd0729020;
                12'd3149: exp <= 22'd0728187;
                12'd3150: exp <= 22'd0727354;
                12'd3151: exp <= 22'd0726521;
                12'd3152: exp <= 22'd0725688;
                12'd3153: exp <= 22'd0724856;
                12'd3154: exp <= 22'd0724023;
                12'd3155: exp <= 22'd0723191;
                12'd3156: exp <= 22'd0722359;
                12'd3157: exp <= 22'd0721527;
                12'd3158: exp <= 22'd0720695;
                12'd3159: exp <= 22'd0719864;
                12'd3160: exp <= 22'd0719032;
                12'd3161: exp <= 22'd0718201;
                12'd3162: exp <= 22'd0717369;
                12'd3163: exp <= 22'd0716538;
                12'd3164: exp <= 22'd0715707;
                12'd3165: exp <= 22'd0714876;
                12'd3166: exp <= 22'd0714046;
                12'd3167: exp <= 22'd0713215;
                12'd3168: exp <= 22'd0712385;
                12'd3169: exp <= 22'd0711555;
                12'd3170: exp <= 22'd0710724;
                12'd3171: exp <= 22'd0709894;
                12'd3172: exp <= 22'd0709065;
                12'd3173: exp <= 22'd0708235;
                12'd3174: exp <= 22'd0707405;
                12'd3175: exp <= 22'd0706576;
                12'd3176: exp <= 22'd0705747;
                12'd3177: exp <= 22'd0704918;
                12'd3178: exp <= 22'd0704089;
                12'd3179: exp <= 22'd0703260;
                12'd3180: exp <= 22'd0702431;
                12'd3181: exp <= 22'd0701602;
                12'd3182: exp <= 22'd0700774;
                12'd3183: exp <= 22'd0699946;
                12'd3184: exp <= 22'd0699117;
                12'd3185: exp <= 22'd0698289;
                12'd3186: exp <= 22'd0697462;
                12'd3187: exp <= 22'd0696634;
                12'd3188: exp <= 22'd0695806;
                12'd3189: exp <= 22'd0694979;
                12'd3190: exp <= 22'd0694151;
                12'd3191: exp <= 22'd0693324;
                12'd3192: exp <= 22'd0692497;
                12'd3193: exp <= 22'd0691670;
                12'd3194: exp <= 22'd0690844;
                12'd3195: exp <= 22'd0690017;
                12'd3196: exp <= 22'd0689190;
                12'd3197: exp <= 22'd0688364;
                12'd3198: exp <= 22'd0687538;
                12'd3199: exp <= 22'd0686712;
                12'd3200: exp <= 22'd0685886;
                12'd3201: exp <= 22'd0685060;
                12'd3202: exp <= 22'd0684234;
                12'd3203: exp <= 22'd0683409;
                12'd3204: exp <= 22'd0682584;
                12'd3205: exp <= 22'd0681758;
                12'd3206: exp <= 22'd0680933;
                12'd3207: exp <= 22'd0680108;
                12'd3208: exp <= 22'd0679284;
                12'd3209: exp <= 22'd0678459;
                12'd3210: exp <= 22'd0677634;
                12'd3211: exp <= 22'd0676810;
                12'd3212: exp <= 22'd0675986;
                12'd3213: exp <= 22'd0675162;
                12'd3214: exp <= 22'd0674338;
                12'd3215: exp <= 22'd0673514;
                12'd3216: exp <= 22'd0672690;
                12'd3217: exp <= 22'd0671867;
                12'd3218: exp <= 22'd0671043;
                12'd3219: exp <= 22'd0670220;
                12'd3220: exp <= 22'd0669397;
                12'd3221: exp <= 22'd0668574;
                12'd3222: exp <= 22'd0667751;
                12'd3223: exp <= 22'd0666928;
                12'd3224: exp <= 22'd0666106;
                12'd3225: exp <= 22'd0665283;
                12'd3226: exp <= 22'd0664461;
                12'd3227: exp <= 22'd0663639;
                12'd3228: exp <= 22'd0662817;
                12'd3229: exp <= 22'd0661995;
                12'd3230: exp <= 22'd0661173;
                12'd3231: exp <= 22'd0660352;
                12'd3232: exp <= 22'd0659530;
                12'd3233: exp <= 22'd0658709;
                12'd3234: exp <= 22'd0657888;
                12'd3235: exp <= 22'd0657067;
                12'd3236: exp <= 22'd0656246;
                12'd3237: exp <= 22'd0655425;
                12'd3238: exp <= 22'd0654604;
                12'd3239: exp <= 22'd0653784;
                12'd3240: exp <= 22'd0652963;
                12'd3241: exp <= 22'd0652143;
                12'd3242: exp <= 22'd0651323;
                12'd3243: exp <= 22'd0650503;
                12'd3244: exp <= 22'd0649683;
                12'd3245: exp <= 22'd0648864;
                12'd3246: exp <= 22'd0648044;
                12'd3247: exp <= 22'd0647225;
                12'd3248: exp <= 22'd0646406;
                12'd3249: exp <= 22'd0645586;
                12'd3250: exp <= 22'd0644768;
                12'd3251: exp <= 22'd0643949;
                12'd3252: exp <= 22'd0643130;
                12'd3253: exp <= 22'd0642311;
                12'd3254: exp <= 22'd0641493;
                12'd3255: exp <= 22'd0640675;
                12'd3256: exp <= 22'd0639857;
                12'd3257: exp <= 22'd0639039;
                12'd3258: exp <= 22'd0638221;
                12'd3259: exp <= 22'd0637403;
                12'd3260: exp <= 22'd0636585;
                12'd3261: exp <= 22'd0635768;
                12'd3262: exp <= 22'd0634951;
                12'd3263: exp <= 22'd0634134;
                12'd3264: exp <= 22'd0633317;
                12'd3265: exp <= 22'd0632500;
                12'd3266: exp <= 22'd0631683;
                12'd3267: exp <= 22'd0630866;
                12'd3268: exp <= 22'd0630050;
                12'd3269: exp <= 22'd0629234;
                12'd3270: exp <= 22'd0628417;
                12'd3271: exp <= 22'd0627601;
                12'd3272: exp <= 22'd0626785;
                12'd3273: exp <= 22'd0625970;
                12'd3274: exp <= 22'd0625154;
                12'd3275: exp <= 22'd0624338;
                12'd3276: exp <= 22'd0623523;
                12'd3277: exp <= 22'd0622708;
                12'd3278: exp <= 22'd0621893;
                12'd3279: exp <= 22'd0621078;
                12'd3280: exp <= 22'd0620263;
                12'd3281: exp <= 22'd0619448;
                12'd3282: exp <= 22'd0618634;
                12'd3283: exp <= 22'd0617819;
                12'd3284: exp <= 22'd0617005;
                12'd3285: exp <= 22'd0616191;
                12'd3286: exp <= 22'd0615377;
                12'd3287: exp <= 22'd0614563;
                12'd3288: exp <= 22'd0613749;
                12'd3289: exp <= 22'd0612936;
                12'd3290: exp <= 22'd0612122;
                12'd3291: exp <= 22'd0611309;
                12'd3292: exp <= 22'd0610496;
                12'd3293: exp <= 22'd0609683;
                12'd3294: exp <= 22'd0608870;
                12'd3295: exp <= 22'd0608057;
                12'd3296: exp <= 22'd0607245;
                12'd3297: exp <= 22'd0606432;
                12'd3298: exp <= 22'd0605620;
                12'd3299: exp <= 22'd0604808;
                12'd3300: exp <= 22'd0603996;
                12'd3301: exp <= 22'd0603184;
                12'd3302: exp <= 22'd0602372;
                12'd3303: exp <= 22'd0601560;
                12'd3304: exp <= 22'd0600749;
                12'd3305: exp <= 22'd0599937;
                12'd3306: exp <= 22'd0599126;
                12'd3307: exp <= 22'd0598315;
                12'd3308: exp <= 22'd0597504;
                12'd3309: exp <= 22'd0596693;
                12'd3310: exp <= 22'd0595882;
                12'd3311: exp <= 22'd0595072;
                12'd3312: exp <= 22'd0594262;
                12'd3313: exp <= 22'd0593451;
                12'd3314: exp <= 22'd0592641;
                12'd3315: exp <= 22'd0591831;
                12'd3316: exp <= 22'd0591021;
                12'd3317: exp <= 22'd0590211;
                12'd3318: exp <= 22'd0589402;
                12'd3319: exp <= 22'd0588592;
                12'd3320: exp <= 22'd0587783;
                12'd3321: exp <= 22'd0586974;
                12'd3322: exp <= 22'd0586165;
                12'd3323: exp <= 22'd0585356;
                12'd3324: exp <= 22'd0584547;
                12'd3325: exp <= 22'd0583739;
                12'd3326: exp <= 22'd0582930;
                12'd3327: exp <= 22'd0582122;
                12'd3328: exp <= 22'd0581314;
                12'd3329: exp <= 22'd0580505;
                12'd3330: exp <= 22'd0579697;
                12'd3331: exp <= 22'd0578890;
                12'd3332: exp <= 22'd0578082;
                12'd3333: exp <= 22'd0577274;
                12'd3334: exp <= 22'd0576467;
                12'd3335: exp <= 22'd0575660;
                12'd3336: exp <= 22'd0574853;
                12'd3337: exp <= 22'd0574046;
                12'd3338: exp <= 22'd0573239;
                12'd3339: exp <= 22'd0572432;
                12'd3340: exp <= 22'd0571625;
                12'd3341: exp <= 22'd0570819;
                12'd3342: exp <= 22'd0570013;
                12'd3343: exp <= 22'd0569207;
                12'd3344: exp <= 22'd0568400;
                12'd3345: exp <= 22'd0567595;
                12'd3346: exp <= 22'd0566789;
                12'd3347: exp <= 22'd0565983;
                12'd3348: exp <= 22'd0565178;
                12'd3349: exp <= 22'd0564372;
                12'd3350: exp <= 22'd0563567;
                12'd3351: exp <= 22'd0562762;
                12'd3352: exp <= 22'd0561957;
                12'd3353: exp <= 22'd0561152;
                12'd3354: exp <= 22'd0560348;
                12'd3355: exp <= 22'd0559543;
                12'd3356: exp <= 22'd0558739;
                12'd3357: exp <= 22'd0557934;
                12'd3358: exp <= 22'd0557130;
                12'd3359: exp <= 22'd0556326;
                12'd3360: exp <= 22'd0555522;
                12'd3361: exp <= 22'd0554719;
                12'd3362: exp <= 22'd0553915;
                12'd3363: exp <= 22'd0553112;
                12'd3364: exp <= 22'd0552308;
                12'd3365: exp <= 22'd0551505;
                12'd3366: exp <= 22'd0550702;
                12'd3367: exp <= 22'd0549899;
                12'd3368: exp <= 22'd0549096;
                12'd3369: exp <= 22'd0548294;
                12'd3370: exp <= 22'd0547491;
                12'd3371: exp <= 22'd0546689;
                12'd3372: exp <= 22'd0545887;
                12'd3373: exp <= 22'd0545085;
                12'd3374: exp <= 22'd0544283;
                12'd3375: exp <= 22'd0543481;
                12'd3376: exp <= 22'd0542679;
                12'd3377: exp <= 22'd0541878;
                12'd3378: exp <= 22'd0541076;
                12'd3379: exp <= 22'd0540275;
                12'd3380: exp <= 22'd0539474;
                12'd3381: exp <= 22'd0538673;
                12'd3382: exp <= 22'd0537872;
                12'd3383: exp <= 22'd0537071;
                12'd3384: exp <= 22'd0536271;
                12'd3385: exp <= 22'd0535470;
                12'd3386: exp <= 22'd0534670;
                12'd3387: exp <= 22'd0533870;
                12'd3388: exp <= 22'd0533069;
                12'd3389: exp <= 22'd0532270;
                12'd3390: exp <= 22'd0531470;
                12'd3391: exp <= 22'd0530670;
                12'd3392: exp <= 22'd0529871;
                12'd3393: exp <= 22'd0529071;
                12'd3394: exp <= 22'd0528272;
                12'd3395: exp <= 22'd0527473;
                12'd3396: exp <= 22'd0526674;
                12'd3397: exp <= 22'd0525875;
                12'd3398: exp <= 22'd0525076;
                12'd3399: exp <= 22'd0524278;
                12'd3400: exp <= 22'd0523479;
                12'd3401: exp <= 22'd0522681;
                12'd3402: exp <= 22'd0521883;
                12'd3403: exp <= 22'd0521085;
                12'd3404: exp <= 22'd0520287;
                12'd3405: exp <= 22'd0519489;
                12'd3406: exp <= 22'd0518692;
                12'd3407: exp <= 22'd0517894;
                12'd3408: exp <= 22'd0517097;
                12'd3409: exp <= 22'd0516299;
                12'd3410: exp <= 22'd0515502;
                12'd3411: exp <= 22'd0514705;
                12'd3412: exp <= 22'd0513909;
                12'd3413: exp <= 22'd0513112;
                12'd3414: exp <= 22'd0512315;
                12'd3415: exp <= 22'd0511519;
                12'd3416: exp <= 22'd0510723;
                12'd3417: exp <= 22'd0509927;
                12'd3418: exp <= 22'd0509131;
                12'd3419: exp <= 22'd0508335;
                12'd3420: exp <= 22'd0507539;
                12'd3421: exp <= 22'd0506743;
                12'd3422: exp <= 22'd0505948;
                12'd3423: exp <= 22'd0505153;
                12'd3424: exp <= 22'd0504357;
                12'd3425: exp <= 22'd0503562;
                12'd3426: exp <= 22'd0502767;
                12'd3427: exp <= 22'd0501973;
                12'd3428: exp <= 22'd0501178;
                12'd3429: exp <= 22'd0500383;
                12'd3430: exp <= 22'd0499589;
                12'd3431: exp <= 22'd0498795;
                12'd3432: exp <= 22'd0498001;
                12'd3433: exp <= 22'd0497207;
                12'd3434: exp <= 22'd0496413;
                12'd3435: exp <= 22'd0495619;
                12'd3436: exp <= 22'd0494825;
                12'd3437: exp <= 22'd0494032;
                12'd3438: exp <= 22'd0493239;
                12'd3439: exp <= 22'd0492445;
                12'd3440: exp <= 22'd0491652;
                12'd3441: exp <= 22'd0490860;
                12'd3442: exp <= 22'd0490067;
                12'd3443: exp <= 22'd0489274;
                12'd3444: exp <= 22'd0488482;
                12'd3445: exp <= 22'd0487689;
                12'd3446: exp <= 22'd0486897;
                12'd3447: exp <= 22'd0486105;
                12'd3448: exp <= 22'd0485313;
                12'd3449: exp <= 22'd0484521;
                12'd3450: exp <= 22'd0483729;
                12'd3451: exp <= 22'd0482938;
                12'd3452: exp <= 22'd0482146;
                12'd3453: exp <= 22'd0481355;
                12'd3454: exp <= 22'd0480564;
                12'd3455: exp <= 22'd0479773;
                12'd3456: exp <= 22'd0478982;
                12'd3457: exp <= 22'd0478191;
                12'd3458: exp <= 22'd0477400;
                12'd3459: exp <= 22'd0476610;
                12'd3460: exp <= 22'd0475820;
                12'd3461: exp <= 22'd0475029;
                12'd3462: exp <= 22'd0474239;
                12'd3463: exp <= 22'd0473449;
                12'd3464: exp <= 22'd0472659;
                12'd3465: exp <= 22'd0471870;
                12'd3466: exp <= 22'd0471080;
                12'd3467: exp <= 22'd0470291;
                12'd3468: exp <= 22'd0469501;
                12'd3469: exp <= 22'd0468712;
                12'd3470: exp <= 22'd0467923;
                12'd3471: exp <= 22'd0467134;
                12'd3472: exp <= 22'd0466346;
                12'd3473: exp <= 22'd0465557;
                12'd3474: exp <= 22'd0464768;
                12'd3475: exp <= 22'd0463980;
                12'd3476: exp <= 22'd0463192;
                12'd3477: exp <= 22'd0462404;
                12'd3478: exp <= 22'd0461616;
                12'd3479: exp <= 22'd0460828;
                12'd3480: exp <= 22'd0460040;
                12'd3481: exp <= 22'd0459253;
                12'd3482: exp <= 22'd0458465;
                12'd3483: exp <= 22'd0457678;
                12'd3484: exp <= 22'd0456891;
                12'd3485: exp <= 22'd0456104;
                12'd3486: exp <= 22'd0455317;
                12'd3487: exp <= 22'd0454530;
                12'd3488: exp <= 22'd0453743;
                12'd3489: exp <= 22'd0452957;
                12'd3490: exp <= 22'd0452171;
                12'd3491: exp <= 22'd0451384;
                12'd3492: exp <= 22'd0450598;
                12'd3493: exp <= 22'd0449812;
                12'd3494: exp <= 22'd0449026;
                12'd3495: exp <= 22'd0448241;
                12'd3496: exp <= 22'd0447455;
                12'd3497: exp <= 22'd0446670;
                12'd3498: exp <= 22'd0445884;
                12'd3499: exp <= 22'd0445099;
                12'd3500: exp <= 22'd0444314;
                12'd3501: exp <= 22'd0443529;
                12'd3502: exp <= 22'd0442745;
                12'd3503: exp <= 22'd0441960;
                12'd3504: exp <= 22'd0441175;
                12'd3505: exp <= 22'd0440391;
                12'd3506: exp <= 22'd0439607;
                12'd3507: exp <= 22'd0438823;
                12'd3508: exp <= 22'd0438039;
                12'd3509: exp <= 22'd0437255;
                12'd3510: exp <= 22'd0436471;
                12'd3511: exp <= 22'd0435688;
                12'd3512: exp <= 22'd0434904;
                12'd3513: exp <= 22'd0434121;
                12'd3514: exp <= 22'd0433338;
                12'd3515: exp <= 22'd0432555;
                12'd3516: exp <= 22'd0431772;
                12'd3517: exp <= 22'd0430989;
                12'd3518: exp <= 22'd0430206;
                12'd3519: exp <= 22'd0429424;
                12'd3520: exp <= 22'd0428641;
                12'd3521: exp <= 22'd0427859;
                12'd3522: exp <= 22'd0427077;
                12'd3523: exp <= 22'd0426295;
                12'd3524: exp <= 22'd0425513;
                12'd3525: exp <= 22'd0424731;
                12'd3526: exp <= 22'd0423950;
                12'd3527: exp <= 22'd0423168;
                12'd3528: exp <= 22'd0422387;
                12'd3529: exp <= 22'd0421606;
                12'd3530: exp <= 22'd0420825;
                12'd3531: exp <= 22'd0420044;
                12'd3532: exp <= 22'd0419263;
                12'd3533: exp <= 22'd0418482;
                12'd3534: exp <= 22'd0417702;
                12'd3535: exp <= 22'd0416921;
                12'd3536: exp <= 22'd0416141;
                12'd3537: exp <= 22'd0415361;
                12'd3538: exp <= 22'd0414581;
                12'd3539: exp <= 22'd0413801;
                12'd3540: exp <= 22'd0413021;
                12'd3541: exp <= 22'd0412242;
                12'd3542: exp <= 22'd0411462;
                12'd3543: exp <= 22'd0410683;
                12'd3544: exp <= 22'd0409904;
                12'd3545: exp <= 22'd0409125;
                12'd3546: exp <= 22'd0408346;
                12'd3547: exp <= 22'd0407567;
                12'd3548: exp <= 22'd0406788;
                12'd3549: exp <= 22'd0406010;
                12'd3550: exp <= 22'd0405231;
                12'd3551: exp <= 22'd0404453;
                12'd3552: exp <= 22'd0403675;
                12'd3553: exp <= 22'd0402897;
                12'd3554: exp <= 22'd0402119;
                12'd3555: exp <= 22'd0401341;
                12'd3556: exp <= 22'd0400563;
                12'd3557: exp <= 22'd0399786;
                12'd3558: exp <= 22'd0399009;
                12'd3559: exp <= 22'd0398231;
                12'd3560: exp <= 22'd0397454;
                12'd3561: exp <= 22'd0396677;
                12'd3562: exp <= 22'd0395900;
                12'd3563: exp <= 22'd0395124;
                12'd3564: exp <= 22'd0394347;
                12'd3565: exp <= 22'd0393571;
                12'd3566: exp <= 22'd0392794;
                12'd3567: exp <= 22'd0392018;
                12'd3568: exp <= 22'd0391242;
                12'd3569: exp <= 22'd0390466;
                12'd3570: exp <= 22'd0389690;
                12'd3571: exp <= 22'd0388915;
                12'd3572: exp <= 22'd0388139;
                12'd3573: exp <= 22'd0387364;
                12'd3574: exp <= 22'd0386588;
                12'd3575: exp <= 22'd0385813;
                12'd3576: exp <= 22'd0385038;
                12'd3577: exp <= 22'd0384263;
                12'd3578: exp <= 22'd0383489;
                12'd3579: exp <= 22'd0382714;
                12'd3580: exp <= 22'd0381940;
                12'd3581: exp <= 22'd0381165;
                12'd3582: exp <= 22'd0380391;
                12'd3583: exp <= 22'd0379617;
                12'd3584: exp <= 22'd0378843;
                12'd3585: exp <= 22'd0378069;
                12'd3586: exp <= 22'd0377295;
                12'd3587: exp <= 22'd0376522;
                12'd3588: exp <= 22'd0375748;
                12'd3589: exp <= 22'd0374975;
                12'd3590: exp <= 22'd0374202;
                12'd3591: exp <= 22'd0373429;
                12'd3592: exp <= 22'd0372656;
                12'd3593: exp <= 22'd0371883;
                12'd3594: exp <= 22'd0371111;
                12'd3595: exp <= 22'd0370338;
                12'd3596: exp <= 22'd0369566;
                12'd3597: exp <= 22'd0368793;
                12'd3598: exp <= 22'd0368021;
                12'd3599: exp <= 22'd0367249;
                12'd3600: exp <= 22'd0366477;
                12'd3601: exp <= 22'd0365706;
                12'd3602: exp <= 22'd0364934;
                12'd3603: exp <= 22'd0364163;
                12'd3604: exp <= 22'd0363391;
                12'd3605: exp <= 22'd0362620;
                12'd3606: exp <= 22'd0361849;
                12'd3607: exp <= 22'd0361078;
                12'd3608: exp <= 22'd0360307;
                12'd3609: exp <= 22'd0359537;
                12'd3610: exp <= 22'd0358766;
                12'd3611: exp <= 22'd0357996;
                12'd3612: exp <= 22'd0357225;
                12'd3613: exp <= 22'd0356455;
                12'd3614: exp <= 22'd0355685;
                12'd3615: exp <= 22'd0354915;
                12'd3616: exp <= 22'd0354145;
                12'd3617: exp <= 22'd0353376;
                12'd3618: exp <= 22'd0352606;
                12'd3619: exp <= 22'd0351837;
                12'd3620: exp <= 22'd0351068;
                12'd3621: exp <= 22'd0350298;
                12'd3622: exp <= 22'd0349529;
                12'd3623: exp <= 22'd0348761;
                12'd3624: exp <= 22'd0347992;
                12'd3625: exp <= 22'd0347223;
                12'd3626: exp <= 22'd0346455;
                12'd3627: exp <= 22'd0345686;
                12'd3628: exp <= 22'd0344918;
                12'd3629: exp <= 22'd0344150;
                12'd3630: exp <= 22'd0343382;
                12'd3631: exp <= 22'd0342614;
                12'd3632: exp <= 22'd0341847;
                12'd3633: exp <= 22'd0341079;
                12'd3634: exp <= 22'd0340312;
                12'd3635: exp <= 22'd0339544;
                12'd3636: exp <= 22'd0338777;
                12'd3637: exp <= 22'd0338010;
                12'd3638: exp <= 22'd0337243;
                12'd3639: exp <= 22'd0336476;
                12'd3640: exp <= 22'd0335710;
                12'd3641: exp <= 22'd0334943;
                12'd3642: exp <= 22'd0334177;
                12'd3643: exp <= 22'd0333411;
                12'd3644: exp <= 22'd0332644;
                12'd3645: exp <= 22'd0331878;
                12'd3646: exp <= 22'd0331112;
                12'd3647: exp <= 22'd0330347;
                12'd3648: exp <= 22'd0329581;
                12'd3649: exp <= 22'd0328816;
                12'd3650: exp <= 22'd0328050;
                12'd3651: exp <= 22'd0327285;
                12'd3652: exp <= 22'd0326520;
                12'd3653: exp <= 22'd0325755;
                12'd3654: exp <= 22'd0324990;
                12'd3655: exp <= 22'd0324225;
                12'd3656: exp <= 22'd0323461;
                12'd3657: exp <= 22'd0322696;
                12'd3658: exp <= 22'd0321932;
                12'd3659: exp <= 22'd0321168;
                12'd3660: exp <= 22'd0320404;
                12'd3661: exp <= 22'd0319640;
                12'd3662: exp <= 22'd0318876;
                12'd3663: exp <= 22'd0318112;
                12'd3664: exp <= 22'd0317349;
                12'd3665: exp <= 22'd0316585;
                12'd3666: exp <= 22'd0315822;
                12'd3667: exp <= 22'd0315059;
                12'd3668: exp <= 22'd0314296;
                12'd3669: exp <= 22'd0313533;
                12'd3670: exp <= 22'd0312770;
                12'd3671: exp <= 22'd0312008;
                12'd3672: exp <= 22'd0311245;
                12'd3673: exp <= 22'd0310483;
                12'd3674: exp <= 22'd0309720;
                12'd3675: exp <= 22'd0308958;
                12'd3676: exp <= 22'd0308196;
                12'd3677: exp <= 22'd0307434;
                12'd3678: exp <= 22'd0306673;
                12'd3679: exp <= 22'd0305911;
                12'd3680: exp <= 22'd0305150;
                12'd3681: exp <= 22'd0304388;
                12'd3682: exp <= 22'd0303627;
                12'd3683: exp <= 22'd0302866;
                12'd3684: exp <= 22'd0302105;
                12'd3685: exp <= 22'd0301344;
                12'd3686: exp <= 22'd0300583;
                12'd3687: exp <= 22'd0299823;
                12'd3688: exp <= 22'd0299062;
                12'd3689: exp <= 22'd0298302;
                12'd3690: exp <= 22'd0297542;
                12'd3691: exp <= 22'd0296782;
                12'd3692: exp <= 22'd0296022;
                12'd3693: exp <= 22'd0295262;
                12'd3694: exp <= 22'd0294502;
                12'd3695: exp <= 22'd0293743;
                12'd3696: exp <= 22'd0292983;
                12'd3697: exp <= 22'd0292224;
                12'd3698: exp <= 22'd0291465;
                12'd3699: exp <= 22'd0290706;
                12'd3700: exp <= 22'd0289947;
                12'd3701: exp <= 22'd0289188;
                12'd3702: exp <= 22'd0288429;
                12'd3703: exp <= 22'd0287671;
                12'd3704: exp <= 22'd0286912;
                12'd3705: exp <= 22'd0286154;
                12'd3706: exp <= 22'd0285396;
                12'd3707: exp <= 22'd0284638;
                12'd3708: exp <= 22'd0283880;
                12'd3709: exp <= 22'd0283122;
                12'd3710: exp <= 22'd0282365;
                12'd3711: exp <= 22'd0281607;
                12'd3712: exp <= 22'd0280850;
                12'd3713: exp <= 22'd0280093;
                12'd3714: exp <= 22'd0279336;
                12'd3715: exp <= 22'd0278579;
                12'd3716: exp <= 22'd0277822;
                12'd3717: exp <= 22'd0277065;
                12'd3718: exp <= 22'd0276308;
                12'd3719: exp <= 22'd0275552;
                12'd3720: exp <= 22'd0274795;
                12'd3721: exp <= 22'd0274039;
                12'd3722: exp <= 22'd0273283;
                12'd3723: exp <= 22'd0272527;
                12'd3724: exp <= 22'd0271771;
                12'd3725: exp <= 22'd0271016;
                12'd3726: exp <= 22'd0270260;
                12'd3727: exp <= 22'd0269505;
                12'd3728: exp <= 22'd0268749;
                12'd3729: exp <= 22'd0267994;
                12'd3730: exp <= 22'd0267239;
                12'd3731: exp <= 22'd0266484;
                12'd3732: exp <= 22'd0265729;
                12'd3733: exp <= 22'd0264975;
                12'd3734: exp <= 22'd0264220;
                12'd3735: exp <= 22'd0263466;
                12'd3736: exp <= 22'd0262711;
                12'd3737: exp <= 22'd0261957;
                12'd3738: exp <= 22'd0261203;
                12'd3739: exp <= 22'd0260449;
                12'd3740: exp <= 22'd0259695;
                12'd3741: exp <= 22'd0258942;
                12'd3742: exp <= 22'd0258188;
                12'd3743: exp <= 22'd0257435;
                12'd3744: exp <= 22'd0256681;
                12'd3745: exp <= 22'd0255928;
                12'd3746: exp <= 22'd0255175;
                12'd3747: exp <= 22'd0254422;
                12'd3748: exp <= 22'd0253670;
                12'd3749: exp <= 22'd0252917;
                12'd3750: exp <= 22'd0252164;
                12'd3751: exp <= 22'd0251412;
                12'd3752: exp <= 22'd0250660;
                12'd3753: exp <= 22'd0249908;
                12'd3754: exp <= 22'd0249156;
                12'd3755: exp <= 22'd0248404;
                12'd3756: exp <= 22'd0247652;
                12'd3757: exp <= 22'd0246900;
                12'd3758: exp <= 22'd0246149;
                12'd3759: exp <= 22'd0245397;
                12'd3760: exp <= 22'd0244646;
                12'd3761: exp <= 22'd0243895;
                12'd3762: exp <= 22'd0243144;
                12'd3763: exp <= 22'd0242393;
                12'd3764: exp <= 22'd0241643;
                12'd3765: exp <= 22'd0240892;
                12'd3766: exp <= 22'd0240141;
                12'd3767: exp <= 22'd0239391;
                12'd3768: exp <= 22'd0238641;
                12'd3769: exp <= 22'd0237891;
                12'd3770: exp <= 22'd0237141;
                12'd3771: exp <= 22'd0236391;
                12'd3772: exp <= 22'd0235641;
                12'd3773: exp <= 22'd0234892;
                12'd3774: exp <= 22'd0234142;
                12'd3775: exp <= 22'd0233393;
                12'd3776: exp <= 22'd0232644;
                12'd3777: exp <= 22'd0231894;
                12'd3778: exp <= 22'd0231146;
                12'd3779: exp <= 22'd0230397;
                12'd3780: exp <= 22'd0229648;
                12'd3781: exp <= 22'd0228899;
                12'd3782: exp <= 22'd0228151;
                12'd3783: exp <= 22'd0227403;
                12'd3784: exp <= 22'd0226654;
                12'd3785: exp <= 22'd0225906;
                12'd3786: exp <= 22'd0225158;
                12'd3787: exp <= 22'd0224411;
                12'd3788: exp <= 22'd0223663;
                12'd3789: exp <= 22'd0222915;
                12'd3790: exp <= 22'd0222168;
                12'd3791: exp <= 22'd0221421;
                12'd3792: exp <= 22'd0220673;
                12'd3793: exp <= 22'd0219926;
                12'd3794: exp <= 22'd0219179;
                12'd3795: exp <= 22'd0218433;
                12'd3796: exp <= 22'd0217686;
                12'd3797: exp <= 22'd0216939;
                12'd3798: exp <= 22'd0216193;
                12'd3799: exp <= 22'd0215447;
                12'd3800: exp <= 22'd0214700;
                12'd3801: exp <= 22'd0213954;
                12'd3802: exp <= 22'd0213208;
                12'd3803: exp <= 22'd0212463;
                12'd3804: exp <= 22'd0211717;
                12'd3805: exp <= 22'd0210971;
                12'd3806: exp <= 22'd0210226;
                12'd3807: exp <= 22'd0209481;
                12'd3808: exp <= 22'd0208736;
                12'd3809: exp <= 22'd0207990;
                12'd3810: exp <= 22'd0207246;
                12'd3811: exp <= 22'd0206501;
                12'd3812: exp <= 22'd0205756;
                12'd3813: exp <= 22'd0205012;
                12'd3814: exp <= 22'd0204267;
                12'd3815: exp <= 22'd0203523;
                12'd3816: exp <= 22'd0202779;
                12'd3817: exp <= 22'd0202035;
                12'd3818: exp <= 22'd0201291;
                12'd3819: exp <= 22'd0200547;
                12'd3820: exp <= 22'd0199803;
                12'd3821: exp <= 22'd0199060;
                12'd3822: exp <= 22'd0198316;
                12'd3823: exp <= 22'd0197573;
                12'd3824: exp <= 22'd0196830;
                12'd3825: exp <= 22'd0196087;
                12'd3826: exp <= 22'd0195344;
                12'd3827: exp <= 22'd0194601;
                12'd3828: exp <= 22'd0193859;
                12'd3829: exp <= 22'd0193116;
                12'd3830: exp <= 22'd0192374;
                12'd3831: exp <= 22'd0191631;
                12'd3832: exp <= 22'd0190889;
                12'd3833: exp <= 22'd0190147;
                12'd3834: exp <= 22'd0189405;
                12'd3835: exp <= 22'd0188664;
                12'd3836: exp <= 22'd0187922;
                12'd3837: exp <= 22'd0187180;
                12'd3838: exp <= 22'd0186439;
                12'd3839: exp <= 22'd0185698;
                12'd3840: exp <= 22'd0184957;
                12'd3841: exp <= 22'd0184216;
                12'd3842: exp <= 22'd0183475;
                12'd3843: exp <= 22'd0182734;
                12'd3844: exp <= 22'd0181993;
                12'd3845: exp <= 22'd0181253;
                12'd3846: exp <= 22'd0180512;
                12'd3847: exp <= 22'd0179772;
                12'd3848: exp <= 22'd0179032;
                12'd3849: exp <= 22'd0178292;
                12'd3850: exp <= 22'd0177552;
                12'd3851: exp <= 22'd0176812;
                12'd3852: exp <= 22'd0176073;
                12'd3853: exp <= 22'd0175333;
                12'd3854: exp <= 22'd0174594;
                12'd3855: exp <= 22'd0173854;
                12'd3856: exp <= 22'd0173115;
                12'd3857: exp <= 22'd0172376;
                12'd3858: exp <= 22'd0171637;
                12'd3859: exp <= 22'd0170899;
                12'd3860: exp <= 22'd0170160;
                12'd3861: exp <= 22'd0169421;
                12'd3862: exp <= 22'd0168683;
                12'd3863: exp <= 22'd0167945;
                12'd3864: exp <= 22'd0167207;
                12'd3865: exp <= 22'd0166469;
                12'd3866: exp <= 22'd0165731;
                12'd3867: exp <= 22'd0164993;
                12'd3868: exp <= 22'd0164255;
                12'd3869: exp <= 22'd0163518;
                12'd3870: exp <= 22'd0162780;
                12'd3871: exp <= 22'd0162043;
                12'd3872: exp <= 22'd0161306;
                12'd3873: exp <= 22'd0160569;
                12'd3874: exp <= 22'd0159832;
                12'd3875: exp <= 22'd0159095;
                12'd3876: exp <= 22'd0158359;
                12'd3877: exp <= 22'd0157622;
                12'd3878: exp <= 22'd0156886;
                12'd3879: exp <= 22'd0156150;
                12'd3880: exp <= 22'd0155413;
                12'd3881: exp <= 22'd0154677;
                12'd3882: exp <= 22'd0153941;
                12'd3883: exp <= 22'd0153206;
                12'd3884: exp <= 22'd0152470;
                12'd3885: exp <= 22'd0151735;
                12'd3886: exp <= 22'd0150999;
                12'd3887: exp <= 22'd0150264;
                12'd3888: exp <= 22'd0149529;
                12'd3889: exp <= 22'd0148794;
                12'd3890: exp <= 22'd0148059;
                12'd3891: exp <= 22'd0147324;
                12'd3892: exp <= 22'd0146589;
                12'd3893: exp <= 22'd0145855;
                12'd3894: exp <= 22'd0145120;
                12'd3895: exp <= 22'd0144386;
                12'd3896: exp <= 22'd0143652;
                12'd3897: exp <= 22'd0142918;
                12'd3898: exp <= 22'd0142184;
                12'd3899: exp <= 22'd0141450;
                12'd3900: exp <= 22'd0140717;
                12'd3901: exp <= 22'd0139983;
                12'd3902: exp <= 22'd0139250;
                12'd3903: exp <= 22'd0138516;
                12'd3904: exp <= 22'd0137783;
                12'd3905: exp <= 22'd0137050;
                12'd3906: exp <= 22'd0136317;
                12'd3907: exp <= 22'd0135584;
                12'd3908: exp <= 22'd0134852;
                12'd3909: exp <= 22'd0134119;
                12'd3910: exp <= 22'd0133387;
                12'd3911: exp <= 22'd0132655;
                12'd3912: exp <= 22'd0131922;
                12'd3913: exp <= 22'd0131190;
                12'd3914: exp <= 22'd0130458;
                12'd3915: exp <= 22'd0129727;
                12'd3916: exp <= 22'd0128995;
                12'd3917: exp <= 22'd0128263;
                12'd3918: exp <= 22'd0127532;
                12'd3919: exp <= 22'd0126801;
                12'd3920: exp <= 22'd0126070;
                12'd3921: exp <= 22'd0125338;
                12'd3922: exp <= 22'd0124608;
                12'd3923: exp <= 22'd0123877;
                12'd3924: exp <= 22'd0123146;
                12'd3925: exp <= 22'd0122415;
                12'd3926: exp <= 22'd0121685;
                12'd3927: exp <= 22'd0120955;
                12'd3928: exp <= 22'd0120225;
                12'd3929: exp <= 22'd0119494;
                12'd3930: exp <= 22'd0118765;
                12'd3931: exp <= 22'd0118035;
                12'd3932: exp <= 22'd0117305;
                12'd3933: exp <= 22'd0116575;
                12'd3934: exp <= 22'd0115846;
                12'd3935: exp <= 22'd0115117;
                12'd3936: exp <= 22'd0114387;
                12'd3937: exp <= 22'd0113658;
                12'd3938: exp <= 22'd0112929;
                12'd3939: exp <= 22'd0112201;
                12'd3940: exp <= 22'd0111472;
                12'd3941: exp <= 22'd0110743;
                12'd3942: exp <= 22'd0110015;
                12'd3943: exp <= 22'd0109286;
                12'd3944: exp <= 22'd0108558;
                12'd3945: exp <= 22'd0107830;
                12'd3946: exp <= 22'd0107102;
                12'd3947: exp <= 22'd0106374;
                12'd3948: exp <= 22'd0105647;
                12'd3949: exp <= 22'd0104919;
                12'd3950: exp <= 22'd0104192;
                12'd3951: exp <= 22'd0103464;
                12'd3952: exp <= 22'd0102737;
                12'd3953: exp <= 22'd0102010;
                12'd3954: exp <= 22'd0101283;
                12'd3955: exp <= 22'd0100556;
                12'd3956: exp <= 22'd0099829;
                12'd3957: exp <= 22'd0099103;
                12'd3958: exp <= 22'd0098376;
                12'd3959: exp <= 22'd0097650;
                12'd3960: exp <= 22'd0096924;
                12'd3961: exp <= 22'd0096197;
                12'd3962: exp <= 22'd0095471;
                12'd3963: exp <= 22'd0094746;
                12'd3964: exp <= 22'd0094020;
                12'd3965: exp <= 22'd0093294;
                12'd3966: exp <= 22'd0092569;
                12'd3967: exp <= 22'd0091843;
                12'd3968: exp <= 22'd0091118;
                12'd3969: exp <= 22'd0090393;
                12'd3970: exp <= 22'd0089668;
                12'd3971: exp <= 22'd0088943;
                12'd3972: exp <= 22'd0088218;
                12'd3973: exp <= 22'd0087494;
                12'd3974: exp <= 22'd0086769;
                12'd3975: exp <= 22'd0086045;
                12'd3976: exp <= 22'd0085320;
                12'd3977: exp <= 22'd0084596;
                12'd3978: exp <= 22'd0083872;
                12'd3979: exp <= 22'd0083148;
                12'd3980: exp <= 22'd0082424;
                12'd3981: exp <= 22'd0081701;
                12'd3982: exp <= 22'd0080977;
                12'd3983: exp <= 22'd0080254;
                12'd3984: exp <= 22'd0079530;
                12'd3985: exp <= 22'd0078807;
                12'd3986: exp <= 22'd0078084;
                12'd3987: exp <= 22'd0077361;
                12'd3988: exp <= 22'd0076639;
                12'd3989: exp <= 22'd0075916;
                12'd3990: exp <= 22'd0075193;
                12'd3991: exp <= 22'd0074471;
                12'd3992: exp <= 22'd0073748;
                12'd3993: exp <= 22'd0073026;
                12'd3994: exp <= 22'd0072304;
                12'd3995: exp <= 22'd0071582;
                12'd3996: exp <= 22'd0070860;
                12'd3997: exp <= 22'd0070139;
                12'd3998: exp <= 22'd0069417;
                12'd3999: exp <= 22'd0068696;
                12'd4000: exp <= 22'd0067974;
                12'd4001: exp <= 22'd0067253;
                12'd4002: exp <= 22'd0066532;
                12'd4003: exp <= 22'd0065811;
                12'd4004: exp <= 22'd0065090;
                12'd4005: exp <= 22'd0064369;
                12'd4006: exp <= 22'd0063649;
                12'd4007: exp <= 22'd0062928;
                12'd4008: exp <= 22'd0062208;
                12'd4009: exp <= 22'd0061488;
                12'd4010: exp <= 22'd0060768;
                12'd4011: exp <= 22'd0060048;
                12'd4012: exp <= 22'd0059328;
                12'd4013: exp <= 22'd0058608;
                12'd4014: exp <= 22'd0057888;
                12'd4015: exp <= 22'd0057169;
                12'd4016: exp <= 22'd0056449;
                12'd4017: exp <= 22'd0055730;
                12'd4018: exp <= 22'd0055011;
                12'd4019: exp <= 22'd0054292;
                12'd4020: exp <= 22'd0053573;
                12'd4021: exp <= 22'd0052854;
                12'd4022: exp <= 22'd0052136;
                12'd4023: exp <= 22'd0051417;
                12'd4024: exp <= 22'd0050699;
                12'd4025: exp <= 22'd0049980;
                12'd4026: exp <= 22'd0049262;
                12'd4027: exp <= 22'd0048544;
                12'd4028: exp <= 22'd0047826;
                12'd4029: exp <= 22'd0047108;
                12'd4030: exp <= 22'd0046391;
                12'd4031: exp <= 22'd0045673;
                12'd4032: exp <= 22'd0044956;
                12'd4033: exp <= 22'd0044238;
                12'd4034: exp <= 22'd0043521;
                12'd4035: exp <= 22'd0042804;
                12'd4036: exp <= 22'd0042087;
                12'd4037: exp <= 22'd0041370;
                12'd4038: exp <= 22'd0040653;
                12'd4039: exp <= 22'd0039937;
                12'd4040: exp <= 22'd0039220;
                12'd4041: exp <= 22'd0038504;
                12'd4042: exp <= 22'd0037788;
                12'd4043: exp <= 22'd0037072;
                12'd4044: exp <= 22'd0036356;
                12'd4045: exp <= 22'd0035640;
                12'd4046: exp <= 22'd0034924;
                12'd4047: exp <= 22'd0034208;
                12'd4048: exp <= 22'd0033493;
                12'd4049: exp <= 22'd0032777;
                12'd4050: exp <= 22'd0032062;
                12'd4051: exp <= 22'd0031347;
                12'd4052: exp <= 22'd0030632;
                12'd4053: exp <= 22'd0029917;
                12'd4054: exp <= 22'd0029202;
                12'd4055: exp <= 22'd0028488;
                12'd4056: exp <= 22'd0027773;
                12'd4057: exp <= 22'd0027059;
                12'd4058: exp <= 22'd0026344;
                12'd4059: exp <= 22'd0025630;
                12'd4060: exp <= 22'd0024916;
                12'd4061: exp <= 22'd0024202;
                12'd4062: exp <= 22'd0023488;
                12'd4063: exp <= 22'd0022775;
                12'd4064: exp <= 22'd0022061;
                12'd4065: exp <= 22'd0021348;
                12'd4066: exp <= 22'd0020634;
                12'd4067: exp <= 22'd0019921;
                12'd4068: exp <= 22'd0019208;
                12'd4069: exp <= 22'd0018495;
                12'd4070: exp <= 22'd0017782;
                12'd4071: exp <= 22'd0017069;
                12'd4072: exp <= 22'd0016357;
                12'd4073: exp <= 22'd0015644;
                12'd4074: exp <= 22'd0014932;
                12'd4075: exp <= 22'd0014220;
                12'd4076: exp <= 22'd0013508;
                12'd4077: exp <= 22'd0012796;
                12'd4078: exp <= 22'd0012084;
                12'd4079: exp <= 22'd0011372;
                12'd4080: exp <= 22'd0010660;
                12'd4081: exp <= 22'd0009949;
                12'd4082: exp <= 22'd0009237;
                12'd4083: exp <= 22'd0008526;
                12'd4084: exp <= 22'd0007815;
                12'd4085: exp <= 22'd0007104;
                12'd4086: exp <= 22'd0006393;
                12'd4087: exp <= 22'd0005682;
                12'd4088: exp <= 22'd0004971;
                12'd4089: exp <= 22'd0004261;
                12'd4090: exp <= 22'd0003550;
                12'd4091: exp <= 22'd0002840;
                12'd4092: exp <= 22'd0002130;
                12'd4093: exp <= 22'd0001420;
                12'd4094: exp <= 22'd0000710;
                12'd4095: exp <= 22'd0000000;
            endcase
        1'b1: //sinexp
            case (addr[19:8])
                12'd0000: exp <= 22'd4194303;
                12'd0001: exp <= 22'd4194302;
                12'd0002: exp <= 22'd4194301;
                12'd0003: exp <= 22'd4194297;
                12'd0004: exp <= 22'd4194293;
                12'd0005: exp <= 22'd4194288;
                12'd0006: exp <= 22'd4194281;
                12'd0007: exp <= 22'd4194273;
                12'd0008: exp <= 22'd4194264;
                12'd0009: exp <= 22'd4194253;
                12'd0010: exp <= 22'd4194241;
                12'd0011: exp <= 22'd4194228;
                12'd0012: exp <= 22'd4194214;
                12'd0013: exp <= 22'd4194199;
                12'd0014: exp <= 22'd4194182;
                12'd0015: exp <= 22'd4194164;
                12'd0016: exp <= 22'd4194145;
                12'd0017: exp <= 22'd4194125;
                12'd0018: exp <= 22'd4194103;
                12'd0019: exp <= 22'd4194080;
                12'd0020: exp <= 22'd4194056;
                12'd0021: exp <= 22'd4194031;
                12'd0022: exp <= 22'd4194004;
                12'd0023: exp <= 22'd4193977;
                12'd0024: exp <= 22'd4193948;
                12'd0025: exp <= 22'd4193917;
                12'd0026: exp <= 22'd4193886;
                12'd0027: exp <= 22'd4193853;
                12'd0028: exp <= 22'd4193819;
                12'd0029: exp <= 22'd4193784;
                12'd0030: exp <= 22'd4193748;
                12'd0031: exp <= 22'd4193710;
                12'd0032: exp <= 22'd4193671;
                12'd0033: exp <= 22'd4193631;
                12'd0034: exp <= 22'd4193590;
                12'd0035: exp <= 22'd4193547;
                12'd0036: exp <= 22'd4193504;
                12'd0037: exp <= 22'd4193459;
                12'd0038: exp <= 22'd4193412;
                12'd0039: exp <= 22'd4193365;
                12'd0040: exp <= 22'd4193316;
                12'd0041: exp <= 22'd4193266;
                12'd0042: exp <= 22'd4193215;
                12'd0043: exp <= 22'd4193163;
                12'd0044: exp <= 22'd4193109;
                12'd0045: exp <= 22'd4193054;
                12'd0046: exp <= 22'd4192998;
                12'd0047: exp <= 22'd4192941;
                12'd0048: exp <= 22'd4192882;
                12'd0049: exp <= 22'd4192822;
                12'd0050: exp <= 22'd4192761;
                12'd0051: exp <= 22'd4192699;
                12'd0052: exp <= 22'd4192635;
                12'd0053: exp <= 22'd4192571;
                12'd0054: exp <= 22'd4192505;
                12'd0055: exp <= 22'd4192437;
                12'd0056: exp <= 22'd4192369;
                12'd0057: exp <= 22'd4192299;
                12'd0058: exp <= 22'd4192228;
                12'd0059: exp <= 22'd4192156;
                12'd0060: exp <= 22'd4192083;
                12'd0061: exp <= 22'd4192008;
                12'd0062: exp <= 22'd4191932;
                12'd0063: exp <= 22'd4191855;
                12'd0064: exp <= 22'd4191777;
                12'd0065: exp <= 22'd4191697;
                12'd0066: exp <= 22'd4191617;
                12'd0067: exp <= 22'd4191535;
                12'd0068: exp <= 22'd4191451;
                12'd0069: exp <= 22'd4191367;
                12'd0070: exp <= 22'd4191281;
                12'd0071: exp <= 22'd4191194;
                12'd0072: exp <= 22'd4191106;
                12'd0073: exp <= 22'd4191017;
                12'd0074: exp <= 22'd4190926;
                12'd0075: exp <= 22'd4190834;
                12'd0076: exp <= 22'd4190741;
                12'd0077: exp <= 22'd4190647;
                12'd0078: exp <= 22'd4190551;
                12'd0079: exp <= 22'd4190454;
                12'd0080: exp <= 22'd4190356;
                12'd0081: exp <= 22'd4190257;
                12'd0082: exp <= 22'd4190157;
                12'd0083: exp <= 22'd4190055;
                12'd0084: exp <= 22'd4189952;
                12'd0085: exp <= 22'd4189848;
                12'd0086: exp <= 22'd4189742;
                12'd0087: exp <= 22'd4189636;
                12'd0088: exp <= 22'd4189528;
                12'd0089: exp <= 22'd4189419;
                12'd0090: exp <= 22'd4189308;
                12'd0091: exp <= 22'd4189197;
                12'd0092: exp <= 22'd4189084;
                12'd0093: exp <= 22'd4188970;
                12'd0094: exp <= 22'd4188855;
                12'd0095: exp <= 22'd4188738;
                12'd0096: exp <= 22'd4188621;
                12'd0097: exp <= 22'd4188502;
                12'd0098: exp <= 22'd4188382;
                12'd0099: exp <= 22'd4188260;
                12'd0100: exp <= 22'd4188138;
                12'd0101: exp <= 22'd4188014;
                12'd0102: exp <= 22'd4187889;
                12'd0103: exp <= 22'd4187762;
                12'd0104: exp <= 22'd4187635;
                12'd0105: exp <= 22'd4187506;
                12'd0106: exp <= 22'd4187376;
                12'd0107: exp <= 22'd4187245;
                12'd0108: exp <= 22'd4187112;
                12'd0109: exp <= 22'd4186978;
                12'd0110: exp <= 22'd4186844;
                12'd0111: exp <= 22'd4186707;
                12'd0112: exp <= 22'd4186570;
                12'd0113: exp <= 22'd4186431;
                12'd0114: exp <= 22'd4186292;
                12'd0115: exp <= 22'd4186150;
                12'd0116: exp <= 22'd4186008;
                12'd0117: exp <= 22'd4185865;
                12'd0118: exp <= 22'd4185720;
                12'd0119: exp <= 22'd4185574;
                12'd0120: exp <= 22'd4185427;
                12'd0121: exp <= 22'd4185278;
                12'd0122: exp <= 22'd4185128;
                12'd0123: exp <= 22'd4184978;
                12'd0124: exp <= 22'd4184825;
                12'd0125: exp <= 22'd4184672;
                12'd0126: exp <= 22'd4184518;
                12'd0127: exp <= 22'd4184362;
                12'd0128: exp <= 22'd4184205;
                12'd0129: exp <= 22'd4184046;
                12'd0130: exp <= 22'd4183887;
                12'd0131: exp <= 22'd4183726;
                12'd0132: exp <= 22'd4183564;
                12'd0133: exp <= 22'd4183401;
                12'd0134: exp <= 22'd4183237;
                12'd0135: exp <= 22'd4183071;
                12'd0136: exp <= 22'd4182904;
                12'd0137: exp <= 22'd4182736;
                12'd0138: exp <= 22'd4182567;
                12'd0139: exp <= 22'd4182396;
                12'd0140: exp <= 22'd4182224;
                12'd0141: exp <= 22'd4182051;
                12'd0142: exp <= 22'd4181877;
                12'd0143: exp <= 22'd4181702;
                12'd0144: exp <= 22'd4181525;
                12'd0145: exp <= 22'd4181347;
                12'd0146: exp <= 22'd4181168;
                12'd0147: exp <= 22'd4180988;
                12'd0148: exp <= 22'd4180806;
                12'd0149: exp <= 22'd4180623;
                12'd0150: exp <= 22'd4180439;
                12'd0151: exp <= 22'd4180254;
                12'd0152: exp <= 22'd4180067;
                12'd0153: exp <= 22'd4179880;
                12'd0154: exp <= 22'd4179691;
                12'd0155: exp <= 22'd4179501;
                12'd0156: exp <= 22'd4179309;
                12'd0157: exp <= 22'd4179117;
                12'd0158: exp <= 22'd4178923;
                12'd0159: exp <= 22'd4178728;
                12'd0160: exp <= 22'd4178531;
                12'd0161: exp <= 22'd4178334;
                12'd0162: exp <= 22'd4178135;
                12'd0163: exp <= 22'd4177935;
                12'd0164: exp <= 22'd4177734;
                12'd0165: exp <= 22'd4177532;
                12'd0166: exp <= 22'd4177328;
                12'd0167: exp <= 22'd4177123;
                12'd0168: exp <= 22'd4176917;
                12'd0169: exp <= 22'd4176710;
                12'd0170: exp <= 22'd4176501;
                12'd0171: exp <= 22'd4176292;
                12'd0172: exp <= 22'd4176081;
                12'd0173: exp <= 22'd4175868;
                12'd0174: exp <= 22'd4175655;
                12'd0175: exp <= 22'd4175440;
                12'd0176: exp <= 22'd4175224;
                12'd0177: exp <= 22'd4175007;
                12'd0178: exp <= 22'd4174789;
                12'd0179: exp <= 22'd4174570;
                12'd0180: exp <= 22'd4174349;
                12'd0181: exp <= 22'd4174127;
                12'd0182: exp <= 22'd4173904;
                12'd0183: exp <= 22'd4173679;
                12'd0184: exp <= 22'd4173454;
                12'd0185: exp <= 22'd4173227;
                12'd0186: exp <= 22'd4172999;
                12'd0187: exp <= 22'd4172769;
                12'd0188: exp <= 22'd4172539;
                12'd0189: exp <= 22'd4172307;
                12'd0190: exp <= 22'd4172074;
                12'd0191: exp <= 22'd4171840;
                12'd0192: exp <= 22'd4171604;
                12'd0193: exp <= 22'd4171368;
                12'd0194: exp <= 22'd4171130;
                12'd0195: exp <= 22'd4170891;
                12'd0196: exp <= 22'd4170651;
                12'd0197: exp <= 22'd4170409;
                12'd0198: exp <= 22'd4170166;
                12'd0199: exp <= 22'd4169922;
                12'd0200: exp <= 22'd4169677;
                12'd0201: exp <= 22'd4169431;
                12'd0202: exp <= 22'd4169183;
                12'd0203: exp <= 22'd4168935;
                12'd0204: exp <= 22'd4168684;
                12'd0205: exp <= 22'd4168433;
                12'd0206: exp <= 22'd4168181;
                12'd0207: exp <= 22'd4167927;
                12'd0208: exp <= 22'd4167672;
                12'd0209: exp <= 22'd4167416;
                12'd0210: exp <= 22'd4167159;
                12'd0211: exp <= 22'd4166900;
                12'd0212: exp <= 22'd4166640;
                12'd0213: exp <= 22'd4166379;
                12'd0214: exp <= 22'd4166117;
                12'd0215: exp <= 22'd4165854;
                12'd0216: exp <= 22'd4165589;
                12'd0217: exp <= 22'd4165323;
                12'd0218: exp <= 22'd4165056;
                12'd0219: exp <= 22'd4164788;
                12'd0220: exp <= 22'd4164518;
                12'd0221: exp <= 22'd4164247;
                12'd0222: exp <= 22'd4163976;
                12'd0223: exp <= 22'd4163702;
                12'd0224: exp <= 22'd4163428;
                12'd0225: exp <= 22'd4163152;
                12'd0226: exp <= 22'd4162876;
                12'd0227: exp <= 22'd4162598;
                12'd0228: exp <= 22'd4162318;
                12'd0229: exp <= 22'd4162038;
                12'd0230: exp <= 22'd4161756;
                12'd0231: exp <= 22'd4161473;
                12'd0232: exp <= 22'd4161189;
                12'd0233: exp <= 22'd4160904;
                12'd0234: exp <= 22'd4160617;
                12'd0235: exp <= 22'd4160330;
                12'd0236: exp <= 22'd4160041;
                12'd0237: exp <= 22'd4159750;
                12'd0238: exp <= 22'd4159459;
                12'd0239: exp <= 22'd4159166;
                12'd0240: exp <= 22'd4158873;
                12'd0241: exp <= 22'd4158578;
                12'd0242: exp <= 22'd4158281;
                12'd0243: exp <= 22'd4157984;
                12'd0244: exp <= 22'd4157685;
                12'd0245: exp <= 22'd4157385;
                12'd0246: exp <= 22'd4157084;
                12'd0247: exp <= 22'd4156782;
                12'd0248: exp <= 22'd4156478;
                12'd0249: exp <= 22'd4156174;
                12'd0250: exp <= 22'd4155868;
                12'd0251: exp <= 22'd4155561;
                12'd0252: exp <= 22'd4155252;
                12'd0253: exp <= 22'd4154943;
                12'd0254: exp <= 22'd4154632;
                12'd0255: exp <= 22'd4154320;
                12'd0256: exp <= 22'd4154007;
                12'd0257: exp <= 22'd4153692;
                12'd0258: exp <= 22'd4153377;
                12'd0259: exp <= 22'd4153060;
                12'd0260: exp <= 22'd4152742;
                12'd0261: exp <= 22'd4152423;
                12'd0262: exp <= 22'd4152102;
                12'd0263: exp <= 22'd4151781;
                12'd0264: exp <= 22'd4151458;
                12'd0265: exp <= 22'd4151134;
                12'd0266: exp <= 22'd4150808;
                12'd0267: exp <= 22'd4150482;
                12'd0268: exp <= 22'd4150154;
                12'd0269: exp <= 22'd4149825;
                12'd0270: exp <= 22'd4149495;
                12'd0271: exp <= 22'd4149164;
                12'd0272: exp <= 22'd4148831;
                12'd0273: exp <= 22'd4148497;
                12'd0274: exp <= 22'd4148163;
                12'd0275: exp <= 22'd4147826;
                12'd0276: exp <= 22'd4147489;
                12'd0277: exp <= 22'd4147150;
                12'd0278: exp <= 22'd4146811;
                12'd0279: exp <= 22'd4146470;
                12'd0280: exp <= 22'd4146128;
                12'd0281: exp <= 22'd4145784;
                12'd0282: exp <= 22'd4145440;
                12'd0283: exp <= 22'd4145094;
                12'd0284: exp <= 22'd4144747;
                12'd0285: exp <= 22'd4144399;
                12'd0286: exp <= 22'd4144049;
                12'd0287: exp <= 22'd4143698;
                12'd0288: exp <= 22'd4143347;
                12'd0289: exp <= 22'd4142994;
                12'd0290: exp <= 22'd4142639;
                12'd0291: exp <= 22'd4142284;
                12'd0292: exp <= 22'd4141927;
                12'd0293: exp <= 22'd4141570;
                12'd0294: exp <= 22'd4141210;
                12'd0295: exp <= 22'd4140850;
                12'd0296: exp <= 22'd4140489;
                12'd0297: exp <= 22'd4140126;
                12'd0298: exp <= 22'd4139762;
                12'd0299: exp <= 22'd4139397;
                12'd0300: exp <= 22'd4139031;
                12'd0301: exp <= 22'd4138664;
                12'd0302: exp <= 22'd4138295;
                12'd0303: exp <= 22'd4137925;
                12'd0304: exp <= 22'd4137554;
                12'd0305: exp <= 22'd4137182;
                12'd0306: exp <= 22'd4136808;
                12'd0307: exp <= 22'd4136434;
                12'd0308: exp <= 22'd4136058;
                12'd0309: exp <= 22'd4135681;
                12'd0310: exp <= 22'd4135302;
                12'd0311: exp <= 22'd4134923;
                12'd0312: exp <= 22'd4134542;
                12'd0313: exp <= 22'd4134160;
                12'd0314: exp <= 22'd4133777;
                12'd0315: exp <= 22'd4133393;
                12'd0316: exp <= 22'd4133008;
                12'd0317: exp <= 22'd4132621;
                12'd0318: exp <= 22'd4132233;
                12'd0319: exp <= 22'd4131844;
                12'd0320: exp <= 22'd4131454;
                12'd0321: exp <= 22'd4131063;
                12'd0322: exp <= 22'd4130670;
                12'd0323: exp <= 22'd4130276;
                12'd0324: exp <= 22'd4129881;
                12'd0325: exp <= 22'd4129485;
                12'd0326: exp <= 22'd4129087;
                12'd0327: exp <= 22'd4128689;
                12'd0328: exp <= 22'd4128289;
                12'd0329: exp <= 22'd4127888;
                12'd0330: exp <= 22'd4127486;
                12'd0331: exp <= 22'd4127082;
                12'd0332: exp <= 22'd4126678;
                12'd0333: exp <= 22'd4126272;
                12'd0334: exp <= 22'd4125865;
                12'd0335: exp <= 22'd4125457;
                12'd0336: exp <= 22'd4125048;
                12'd0337: exp <= 22'd4124637;
                12'd0338: exp <= 22'd4124225;
                12'd0339: exp <= 22'd4123812;
                12'd0340: exp <= 22'd4123398;
                12'd0341: exp <= 22'd4122983;
                12'd0342: exp <= 22'd4122566;
                12'd0343: exp <= 22'd4122149;
                12'd0344: exp <= 22'd4121730;
                12'd0345: exp <= 22'd4121310;
                12'd0346: exp <= 22'd4120889;
                12'd0347: exp <= 22'd4120466;
                12'd0348: exp <= 22'd4120042;
                12'd0349: exp <= 22'd4119618;
                12'd0350: exp <= 22'd4119192;
                12'd0351: exp <= 22'd4118764;
                12'd0352: exp <= 22'd4118336;
                12'd0353: exp <= 22'd4117906;
                12'd0354: exp <= 22'd4117476;
                12'd0355: exp <= 22'd4117044;
                12'd0356: exp <= 22'd4116610;
                12'd0357: exp <= 22'd4116176;
                12'd0358: exp <= 22'd4115740;
                12'd0359: exp <= 22'd4115304;
                12'd0360: exp <= 22'd4114866;
                12'd0361: exp <= 22'd4114427;
                12'd0362: exp <= 22'd4113986;
                12'd0363: exp <= 22'd4113545;
                12'd0364: exp <= 22'd4113102;
                12'd0365: exp <= 22'd4112658;
                12'd0366: exp <= 22'd4112213;
                12'd0367: exp <= 22'd4111767;
                12'd0368: exp <= 22'd4111320;
                12'd0369: exp <= 22'd4110871;
                12'd0370: exp <= 22'd4110421;
                12'd0371: exp <= 22'd4109970;
                12'd0372: exp <= 22'd4109518;
                12'd0373: exp <= 22'd4109065;
                12'd0374: exp <= 22'd4108610;
                12'd0375: exp <= 22'd4108155;
                12'd0376: exp <= 22'd4107698;
                12'd0377: exp <= 22'd4107240;
                12'd0378: exp <= 22'd4106781;
                12'd0379: exp <= 22'd4106320;
                12'd0380: exp <= 22'd4105859;
                12'd0381: exp <= 22'd4105396;
                12'd0382: exp <= 22'd4104932;
                12'd0383: exp <= 22'd4104467;
                12'd0384: exp <= 22'd4104000;
                12'd0385: exp <= 22'd4103533;
                12'd0386: exp <= 22'd4103064;
                12'd0387: exp <= 22'd4102594;
                12'd0388: exp <= 22'd4102123;
                12'd0389: exp <= 22'd4101651;
                12'd0390: exp <= 22'd4101178;
                12'd0391: exp <= 22'd4100703;
                12'd0392: exp <= 22'd4100227;
                12'd0393: exp <= 22'd4099750;
                12'd0394: exp <= 22'd4099272;
                12'd0395: exp <= 22'd4098793;
                12'd0396: exp <= 22'd4098312;
                12'd0397: exp <= 22'd4097831;
                12'd0398: exp <= 22'd4097348;
                12'd0399: exp <= 22'd4096864;
                12'd0400: exp <= 22'd4096379;
                12'd0401: exp <= 22'd4095892;
                12'd0402: exp <= 22'd4095405;
                12'd0403: exp <= 22'd4094916;
                12'd0404: exp <= 22'd4094426;
                12'd0405: exp <= 22'd4093935;
                12'd0406: exp <= 22'd4093443;
                12'd0407: exp <= 22'd4092949;
                12'd0408: exp <= 22'd4092455;
                12'd0409: exp <= 22'd4091959;
                12'd0410: exp <= 22'd4091462;
                12'd0411: exp <= 22'd4090964;
                12'd0412: exp <= 22'd4090465;
                12'd0413: exp <= 22'd4089964;
                12'd0414: exp <= 22'd4089463;
                12'd0415: exp <= 22'd4088960;
                12'd0416: exp <= 22'd4088456;
                12'd0417: exp <= 22'd4087951;
                12'd0418: exp <= 22'd4087444;
                12'd0419: exp <= 22'd4086937;
                12'd0420: exp <= 22'd4086428;
                12'd0421: exp <= 22'd4085919;
                12'd0422: exp <= 22'd4085408;
                12'd0423: exp <= 22'd4084895;
                12'd0424: exp <= 22'd4084382;
                12'd0425: exp <= 22'd4083868;
                12'd0426: exp <= 22'd4083352;
                12'd0427: exp <= 22'd4082835;
                12'd0428: exp <= 22'd4082317;
                12'd0429: exp <= 22'd4081798;
                12'd0430: exp <= 22'd4081277;
                12'd0431: exp <= 22'd4080756;
                12'd0432: exp <= 22'd4080233;
                12'd0433: exp <= 22'd4079709;
                12'd0434: exp <= 22'd4079184;
                12'd0435: exp <= 22'd4078658;
                12'd0436: exp <= 22'd4078131;
                12'd0437: exp <= 22'd4077602;
                12'd0438: exp <= 22'd4077073;
                12'd0439: exp <= 22'd4076542;
                12'd0440: exp <= 22'd4076010;
                12'd0441: exp <= 22'd4075477;
                12'd0442: exp <= 22'd4074942;
                12'd0443: exp <= 22'd4074407;
                12'd0444: exp <= 22'd4073870;
                12'd0445: exp <= 22'd4073332;
                12'd0446: exp <= 22'd4072793;
                12'd0447: exp <= 22'd4072253;
                12'd0448: exp <= 22'd4071712;
                12'd0449: exp <= 22'd4071170;
                12'd0450: exp <= 22'd4070626;
                12'd0451: exp <= 22'd4070081;
                12'd0452: exp <= 22'd4069535;
                12'd0453: exp <= 22'd4068988;
                12'd0454: exp <= 22'd4068440;
                12'd0455: exp <= 22'd4067890;
                12'd0456: exp <= 22'd4067340;
                12'd0457: exp <= 22'd4066788;
                12'd0458: exp <= 22'd4066235;
                12'd0459: exp <= 22'd4065681;
                12'd0460: exp <= 22'd4065126;
                12'd0461: exp <= 22'd4064569;
                12'd0462: exp <= 22'd4064012;
                12'd0463: exp <= 22'd4063453;
                12'd0464: exp <= 22'd4062893;
                12'd0465: exp <= 22'd4062332;
                12'd0466: exp <= 22'd4061770;
                12'd0467: exp <= 22'd4061207;
                12'd0468: exp <= 22'd4060642;
                12'd0469: exp <= 22'd4060077;
                12'd0470: exp <= 22'd4059510;
                12'd0471: exp <= 22'd4058942;
                12'd0472: exp <= 22'd4058373;
                12'd0473: exp <= 22'd4057803;
                12'd0474: exp <= 22'd4057231;
                12'd0475: exp <= 22'd4056659;
                12'd0476: exp <= 22'd4056085;
                12'd0477: exp <= 22'd4055510;
                12'd0478: exp <= 22'd4054934;
                12'd0479: exp <= 22'd4054357;
                12'd0480: exp <= 22'd4053779;
                12'd0481: exp <= 22'd4053199;
                12'd0482: exp <= 22'd4052619;
                12'd0483: exp <= 22'd4052037;
                12'd0484: exp <= 22'd4051454;
                12'd0485: exp <= 22'd4050870;
                12'd0486: exp <= 22'd4050285;
                12'd0487: exp <= 22'd4049698;
                12'd0488: exp <= 22'd4049111;
                12'd0489: exp <= 22'd4048522;
                12'd0490: exp <= 22'd4047932;
                12'd0491: exp <= 22'd4047341;
                12'd0492: exp <= 22'd4046749;
                12'd0493: exp <= 22'd4046156;
                12'd0494: exp <= 22'd4045562;
                12'd0495: exp <= 22'd4044966;
                12'd0496: exp <= 22'd4044369;
                12'd0497: exp <= 22'd4043772;
                12'd0498: exp <= 22'd4043173;
                12'd0499: exp <= 22'd4042572;
                12'd0500: exp <= 22'd4041971;
                12'd0501: exp <= 22'd4041369;
                12'd0502: exp <= 22'd4040765;
                12'd0503: exp <= 22'd4040161;
                12'd0504: exp <= 22'd4039555;
                12'd0505: exp <= 22'd4038948;
                12'd0506: exp <= 22'd4038340;
                12'd0507: exp <= 22'd4037730;
                12'd0508: exp <= 22'd4037120;
                12'd0509: exp <= 22'd4036508;
                12'd0510: exp <= 22'd4035896;
                12'd0511: exp <= 22'd4035282;
                12'd0512: exp <= 22'd4034667;
                12'd0513: exp <= 22'd4034051;
                12'd0514: exp <= 22'd4033433;
                12'd0515: exp <= 22'd4032815;
                12'd0516: exp <= 22'd4032196;
                12'd0517: exp <= 22'd4031575;
                12'd0518: exp <= 22'd4030953;
                12'd0519: exp <= 22'd4030330;
                12'd0520: exp <= 22'd4029706;
                12'd0521: exp <= 22'd4029081;
                12'd0522: exp <= 22'd4028454;
                12'd0523: exp <= 22'd4027827;
                12'd0524: exp <= 22'd4027198;
                12'd0525: exp <= 22'd4026569;
                12'd0526: exp <= 22'd4025938;
                12'd0527: exp <= 22'd4025306;
                12'd0528: exp <= 22'd4024672;
                12'd0529: exp <= 22'd4024038;
                12'd0530: exp <= 22'd4023403;
                12'd0531: exp <= 22'd4022766;
                12'd0532: exp <= 22'd4022128;
                12'd0533: exp <= 22'd4021490;
                12'd0534: exp <= 22'd4020850;
                12'd0535: exp <= 22'd4020209;
                12'd0536: exp <= 22'd4019566;
                12'd0537: exp <= 22'd4018923;
                12'd0538: exp <= 22'd4018278;
                12'd0539: exp <= 22'd4017633;
                12'd0540: exp <= 22'd4016986;
                12'd0541: exp <= 22'd4016338;
                12'd0542: exp <= 22'd4015689;
                12'd0543: exp <= 22'd4015039;
                12'd0544: exp <= 22'd4014388;
                12'd0545: exp <= 22'd4013735;
                12'd0546: exp <= 22'd4013082;
                12'd0547: exp <= 22'd4012427;
                12'd0548: exp <= 22'd4011771;
                12'd0549: exp <= 22'd4011115;
                12'd0550: exp <= 22'd4010457;
                12'd0551: exp <= 22'd4009797;
                12'd0552: exp <= 22'd4009137;
                12'd0553: exp <= 22'd4008476;
                12'd0554: exp <= 22'd4007813;
                12'd0555: exp <= 22'd4007150;
                12'd0556: exp <= 22'd4006485;
                12'd0557: exp <= 22'd4005819;
                12'd0558: exp <= 22'd4005152;
                12'd0559: exp <= 22'd4004484;
                12'd0560: exp <= 22'd4003814;
                12'd0561: exp <= 22'd4003144;
                12'd0562: exp <= 22'd4002473;
                12'd0563: exp <= 22'd4001800;
                12'd0564: exp <= 22'd4001126;
                12'd0565: exp <= 22'd4000451;
                12'd0566: exp <= 22'd3999775;
                12'd0567: exp <= 22'd3999098;
                12'd0568: exp <= 22'd3998420;
                12'd0569: exp <= 22'd3997741;
                12'd0570: exp <= 22'd3997060;
                12'd0571: exp <= 22'd3996379;
                12'd0572: exp <= 22'd3995696;
                12'd0573: exp <= 22'd3995012;
                12'd0574: exp <= 22'd3994327;
                12'd0575: exp <= 22'd3993641;
                12'd0576: exp <= 22'd3992954;
                12'd0577: exp <= 22'd3992266;
                12'd0578: exp <= 22'd3991576;
                12'd0579: exp <= 22'd3990886;
                12'd0580: exp <= 22'd3990194;
                12'd0581: exp <= 22'd3989501;
                12'd0582: exp <= 22'd3988808;
                12'd0583: exp <= 22'd3988113;
                12'd0584: exp <= 22'd3987417;
                12'd0585: exp <= 22'd3986719;
                12'd0586: exp <= 22'd3986021;
                12'd0587: exp <= 22'd3985322;
                12'd0588: exp <= 22'd3984621;
                12'd0589: exp <= 22'd3983919;
                12'd0590: exp <= 22'd3983217;
                12'd0591: exp <= 22'd3982513;
                12'd0592: exp <= 22'd3981808;
                12'd0593: exp <= 22'd3981102;
                12'd0594: exp <= 22'd3980395;
                12'd0595: exp <= 22'd3979686;
                12'd0596: exp <= 22'd3978977;
                12'd0597: exp <= 22'd3978267;
                12'd0598: exp <= 22'd3977555;
                12'd0599: exp <= 22'd3976842;
                12'd0600: exp <= 22'd3976128;
                12'd0601: exp <= 22'd3975413;
                12'd0602: exp <= 22'd3974697;
                12'd0603: exp <= 22'd3973980;
                12'd0604: exp <= 22'd3973262;
                12'd0605: exp <= 22'd3972543;
                12'd0606: exp <= 22'd3971822;
                12'd0607: exp <= 22'd3971101;
                12'd0608: exp <= 22'd3970378;
                12'd0609: exp <= 22'd3969654;
                12'd0610: exp <= 22'd3968930;
                12'd0611: exp <= 22'd3968204;
                12'd0612: exp <= 22'd3967477;
                12'd0613: exp <= 22'd3966748;
                12'd0614: exp <= 22'd3966019;
                12'd0615: exp <= 22'd3965289;
                12'd0616: exp <= 22'd3964557;
                12'd0617: exp <= 22'd3963825;
                12'd0618: exp <= 22'd3963091;
                12'd0619: exp <= 22'd3962356;
                12'd0620: exp <= 22'd3961621;
                12'd0621: exp <= 22'd3960884;
                12'd0622: exp <= 22'd3960146;
                12'd0623: exp <= 22'd3959406;
                12'd0624: exp <= 22'd3958666;
                12'd0625: exp <= 22'd3957925;
                12'd0626: exp <= 22'd3957182;
                12'd0627: exp <= 22'd3956439;
                12'd0628: exp <= 22'd3955694;
                12'd0629: exp <= 22'd3954949;
                12'd0630: exp <= 22'd3954202;
                12'd0631: exp <= 22'd3953454;
                12'd0632: exp <= 22'd3952705;
                12'd0633: exp <= 22'd3951955;
                12'd0634: exp <= 22'd3951204;
                12'd0635: exp <= 22'd3950452;
                12'd0636: exp <= 22'd3949698;
                12'd0637: exp <= 22'd3948944;
                12'd0638: exp <= 22'd3948188;
                12'd0639: exp <= 22'd3947432;
                12'd0640: exp <= 22'd3946674;
                12'd0641: exp <= 22'd3945915;
                12'd0642: exp <= 22'd3945155;
                12'd0643: exp <= 22'd3944394;
                12'd0644: exp <= 22'd3943632;
                12'd0645: exp <= 22'd3942869;
                12'd0646: exp <= 22'd3942105;
                12'd0647: exp <= 22'd3941340;
                12'd0648: exp <= 22'd3940573;
                12'd0649: exp <= 22'd3939806;
                12'd0650: exp <= 22'd3939037;
                12'd0651: exp <= 22'd3938268;
                12'd0652: exp <= 22'd3937497;
                12'd0653: exp <= 22'd3936725;
                12'd0654: exp <= 22'd3935952;
                12'd0655: exp <= 22'd3935178;
                12'd0656: exp <= 22'd3934403;
                12'd0657: exp <= 22'd3933627;
                12'd0658: exp <= 22'd3932850;
                12'd0659: exp <= 22'd3932072;
                12'd0660: exp <= 22'd3931292;
                12'd0661: exp <= 22'd3930512;
                12'd0662: exp <= 22'd3929730;
                12'd0663: exp <= 22'd3928948;
                12'd0664: exp <= 22'd3928164;
                12'd0665: exp <= 22'd3927379;
                12'd0666: exp <= 22'd3926593;
                12'd0667: exp <= 22'd3925806;
                12'd0668: exp <= 22'd3925018;
                12'd0669: exp <= 22'd3924229;
                12'd0670: exp <= 22'd3923439;
                12'd0671: exp <= 22'd3922648;
                12'd0672: exp <= 22'd3921856;
                12'd0673: exp <= 22'd3921062;
                12'd0674: exp <= 22'd3920268;
                12'd0675: exp <= 22'd3919472;
                12'd0676: exp <= 22'd3918676;
                12'd0677: exp <= 22'd3917878;
                12'd0678: exp <= 22'd3917079;
                12'd0679: exp <= 22'd3916280;
                12'd0680: exp <= 22'd3915479;
                12'd0681: exp <= 22'd3914677;
                12'd0682: exp <= 22'd3913874;
                12'd0683: exp <= 22'd3913070;
                12'd0684: exp <= 22'd3912265;
                12'd0685: exp <= 22'd3911458;
                12'd0686: exp <= 22'd3910651;
                12'd0687: exp <= 22'd3909843;
                12'd0688: exp <= 22'd3909033;
                12'd0689: exp <= 22'd3908223;
                12'd0690: exp <= 22'd3907411;
                12'd0691: exp <= 22'd3906599;
                12'd0692: exp <= 22'd3905785;
                12'd0693: exp <= 22'd3904970;
                12'd0694: exp <= 22'd3904155;
                12'd0695: exp <= 22'd3903338;
                12'd0696: exp <= 22'd3902520;
                12'd0697: exp <= 22'd3901701;
                12'd0698: exp <= 22'd3900881;
                12'd0699: exp <= 22'd3900060;
                12'd0700: exp <= 22'd3899238;
                12'd0701: exp <= 22'd3898414;
                12'd0702: exp <= 22'd3897590;
                12'd0703: exp <= 22'd3896765;
                12'd0704: exp <= 22'd3895938;
                12'd0705: exp <= 22'd3895111;
                12'd0706: exp <= 22'd3894282;
                12'd0707: exp <= 22'd3893453;
                12'd0708: exp <= 22'd3892622;
                12'd0709: exp <= 22'd3891790;
                12'd0710: exp <= 22'd3890958;
                12'd0711: exp <= 22'd3890124;
                12'd0712: exp <= 22'd3889289;
                12'd0713: exp <= 22'd3888453;
                12'd0714: exp <= 22'd3887616;
                12'd0715: exp <= 22'd3886778;
                12'd0716: exp <= 22'd3885939;
                12'd0717: exp <= 22'd3885099;
                12'd0718: exp <= 22'd3884258;
                12'd0719: exp <= 22'd3883416;
                12'd0720: exp <= 22'd3882572;
                12'd0721: exp <= 22'd3881728;
                12'd0722: exp <= 22'd3880883;
                12'd0723: exp <= 22'd3880036;
                12'd0724: exp <= 22'd3879189;
                12'd0725: exp <= 22'd3878340;
                12'd0726: exp <= 22'd3877491;
                12'd0727: exp <= 22'd3876640;
                12'd0728: exp <= 22'd3875788;
                12'd0729: exp <= 22'd3874936;
                12'd0730: exp <= 22'd3874082;
                12'd0731: exp <= 22'd3873227;
                12'd0732: exp <= 22'd3872371;
                12'd0733: exp <= 22'd3871514;
                12'd0734: exp <= 22'd3870656;
                12'd0735: exp <= 22'd3869797;
                12'd0736: exp <= 22'd3868937;
                12'd0737: exp <= 22'd3868076;
                12'd0738: exp <= 22'd3867214;
                12'd0739: exp <= 22'd3866351;
                12'd0740: exp <= 22'd3865487;
                12'd0741: exp <= 22'd3864622;
                12'd0742: exp <= 22'd3863755;
                12'd0743: exp <= 22'd3862888;
                12'd0744: exp <= 22'd3862020;
                12'd0745: exp <= 22'd3861150;
                12'd0746: exp <= 22'd3860280;
                12'd0747: exp <= 22'd3859408;
                12'd0748: exp <= 22'd3858536;
                12'd0749: exp <= 22'd3857662;
                12'd0750: exp <= 22'd3856788;
                12'd0751: exp <= 22'd3855912;
                12'd0752: exp <= 22'd3855036;
                12'd0753: exp <= 22'd3854158;
                12'd0754: exp <= 22'd3853279;
                12'd0755: exp <= 22'd3852400;
                12'd0756: exp <= 22'd3851519;
                12'd0757: exp <= 22'd3850637;
                12'd0758: exp <= 22'd3849754;
                12'd0759: exp <= 22'd3848870;
                12'd0760: exp <= 22'd3847985;
                12'd0761: exp <= 22'd3847099;
                12'd0762: exp <= 22'd3846212;
                12'd0763: exp <= 22'd3845324;
                12'd0764: exp <= 22'd3844435;
                12'd0765: exp <= 22'd3843545;
                12'd0766: exp <= 22'd3842654;
                12'd0767: exp <= 22'd3841762;
                12'd0768: exp <= 22'd3840869;
                12'd0769: exp <= 22'd3839975;
                12'd0770: exp <= 22'd3839080;
                12'd0771: exp <= 22'd3838184;
                12'd0772: exp <= 22'd3837286;
                12'd0773: exp <= 22'd3836388;
                12'd0774: exp <= 22'd3835489;
                12'd0775: exp <= 22'd3834589;
                12'd0776: exp <= 22'd3833687;
                12'd0777: exp <= 22'd3832785;
                12'd0778: exp <= 22'd3831882;
                12'd0779: exp <= 22'd3830977;
                12'd0780: exp <= 22'd3830072;
                12'd0781: exp <= 22'd3829165;
                12'd0782: exp <= 22'd3828258;
                12'd0783: exp <= 22'd3827350;
                12'd0784: exp <= 22'd3826440;
                12'd0785: exp <= 22'd3825530;
                12'd0786: exp <= 22'd3824618;
                12'd0787: exp <= 22'd3823706;
                12'd0788: exp <= 22'd3822792;
                12'd0789: exp <= 22'd3821878;
                12'd0790: exp <= 22'd3820962;
                12'd0791: exp <= 22'd3820045;
                12'd0792: exp <= 22'd3819128;
                12'd0793: exp <= 22'd3818209;
                12'd0794: exp <= 22'd3817290;
                12'd0795: exp <= 22'd3816369;
                12'd0796: exp <= 22'd3815447;
                12'd0797: exp <= 22'd3814525;
                12'd0798: exp <= 22'd3813601;
                12'd0799: exp <= 22'd3812676;
                12'd0800: exp <= 22'd3811751;
                12'd0801: exp <= 22'd3810824;
                12'd0802: exp <= 22'd3809896;
                12'd0803: exp <= 22'd3808968;
                12'd0804: exp <= 22'd3808038;
                12'd0805: exp <= 22'd3807107;
                12'd0806: exp <= 22'd3806175;
                12'd0807: exp <= 22'd3805243;
                12'd0808: exp <= 22'd3804309;
                12'd0809: exp <= 22'd3803374;
                12'd0810: exp <= 22'd3802438;
                12'd0811: exp <= 22'd3801502;
                12'd0812: exp <= 22'd3800564;
                12'd0813: exp <= 22'd3799625;
                12'd0814: exp <= 22'd3798685;
                12'd0815: exp <= 22'd3797745;
                12'd0816: exp <= 22'd3796803;
                12'd0817: exp <= 22'd3795860;
                12'd0818: exp <= 22'd3794916;
                12'd0819: exp <= 22'd3793972;
                12'd0820: exp <= 22'd3793026;
                12'd0821: exp <= 22'd3792079;
                12'd0822: exp <= 22'd3791131;
                12'd0823: exp <= 22'd3790183;
                12'd0824: exp <= 22'd3789233;
                12'd0825: exp <= 22'd3788282;
                12'd0826: exp <= 22'd3787331;
                12'd0827: exp <= 22'd3786378;
                12'd0828: exp <= 22'd3785424;
                12'd0829: exp <= 22'd3784469;
                12'd0830: exp <= 22'd3783514;
                12'd0831: exp <= 22'd3782557;
                12'd0832: exp <= 22'd3781599;
                12'd0833: exp <= 22'd3780641;
                12'd0834: exp <= 22'd3779681;
                12'd0835: exp <= 22'd3778720;
                12'd0836: exp <= 22'd3777759;
                12'd0837: exp <= 22'd3776796;
                12'd0838: exp <= 22'd3775832;
                12'd0839: exp <= 22'd3774868;
                12'd0840: exp <= 22'd3773902;
                12'd0841: exp <= 22'd3772936;
                12'd0842: exp <= 22'd3771968;
                12'd0843: exp <= 22'd3770999;
                12'd0844: exp <= 22'd3770030;
                12'd0845: exp <= 22'd3769059;
                12'd0846: exp <= 22'd3768088;
                12'd0847: exp <= 22'd3767115;
                12'd0848: exp <= 22'd3766142;
                12'd0849: exp <= 22'd3765168;
                12'd0850: exp <= 22'd3764192;
                12'd0851: exp <= 22'd3763216;
                12'd0852: exp <= 22'd3762238;
                12'd0853: exp <= 22'd3761260;
                12'd0854: exp <= 22'd3760281;
                12'd0855: exp <= 22'd3759300;
                12'd0856: exp <= 22'd3758319;
                12'd0857: exp <= 22'd3757337;
                12'd0858: exp <= 22'd3756353;
                12'd0859: exp <= 22'd3755369;
                12'd0860: exp <= 22'd3754384;
                12'd0861: exp <= 22'd3753398;
                12'd0862: exp <= 22'd3752411;
                12'd0863: exp <= 22'd3751422;
                12'd0864: exp <= 22'd3750433;
                12'd0865: exp <= 22'd3749443;
                12'd0866: exp <= 22'd3748452;
                12'd0867: exp <= 22'd3747460;
                12'd0868: exp <= 22'd3746467;
                12'd0869: exp <= 22'd3745473;
                12'd0870: exp <= 22'd3744478;
                12'd0871: exp <= 22'd3743482;
                12'd0872: exp <= 22'd3742485;
                12'd0873: exp <= 22'd3741488;
                12'd0874: exp <= 22'd3740489;
                12'd0875: exp <= 22'd3739489;
                12'd0876: exp <= 22'd3738488;
                12'd0877: exp <= 22'd3737487;
                12'd0878: exp <= 22'd3736484;
                12'd0879: exp <= 22'd3735480;
                12'd0880: exp <= 22'd3734476;
                12'd0881: exp <= 22'd3733470;
                12'd0882: exp <= 22'd3732464;
                12'd0883: exp <= 22'd3731456;
                12'd0884: exp <= 22'd3730448;
                12'd0885: exp <= 22'd3729438;
                12'd0886: exp <= 22'd3728428;
                12'd0887: exp <= 22'd3727416;
                12'd0888: exp <= 22'd3726404;
                12'd0889: exp <= 22'd3725391;
                12'd0890: exp <= 22'd3724377;
                12'd0891: exp <= 22'd3723362;
                12'd0892: exp <= 22'd3722345;
                12'd0893: exp <= 22'd3721328;
                12'd0894: exp <= 22'd3720310;
                12'd0895: exp <= 22'd3719291;
                12'd0896: exp <= 22'd3718271;
                12'd0897: exp <= 22'd3717251;
                12'd0898: exp <= 22'd3716229;
                12'd0899: exp <= 22'd3715206;
                12'd0900: exp <= 22'd3714182;
                12'd0901: exp <= 22'd3713157;
                12'd0902: exp <= 22'd3712132;
                12'd0903: exp <= 22'd3711105;
                12'd0904: exp <= 22'd3710078;
                12'd0905: exp <= 22'd3709049;
                12'd0906: exp <= 22'd3708020;
                12'd0907: exp <= 22'd3706989;
                12'd0908: exp <= 22'd3705958;
                12'd0909: exp <= 22'd3704926;
                12'd0910: exp <= 22'd3703892;
                12'd0911: exp <= 22'd3702858;
                12'd0912: exp <= 22'd3701823;
                12'd0913: exp <= 22'd3700787;
                12'd0914: exp <= 22'd3699750;
                12'd0915: exp <= 22'd3698712;
                12'd0916: exp <= 22'd3697673;
                12'd0917: exp <= 22'd3696633;
                12'd0918: exp <= 22'd3695592;
                12'd0919: exp <= 22'd3694551;
                12'd0920: exp <= 22'd3693508;
                12'd0921: exp <= 22'd3692465;
                12'd0922: exp <= 22'd3691420;
                12'd0923: exp <= 22'd3690374;
                12'd0924: exp <= 22'd3689328;
                12'd0925: exp <= 22'd3688281;
                12'd0926: exp <= 22'd3687232;
                12'd0927: exp <= 22'd3686183;
                12'd0928: exp <= 22'd3685133;
                12'd0929: exp <= 22'd3684082;
                12'd0930: exp <= 22'd3683030;
                12'd0931: exp <= 22'd3681977;
                12'd0932: exp <= 22'd3680923;
                12'd0933: exp <= 22'd3679868;
                12'd0934: exp <= 22'd3678813;
                12'd0935: exp <= 22'd3677756;
                12'd0936: exp <= 22'd3676698;
                12'd0937: exp <= 22'd3675640;
                12'd0938: exp <= 22'd3674580;
                12'd0939: exp <= 22'd3673520;
                12'd0940: exp <= 22'd3672458;
                12'd0941: exp <= 22'd3671396;
                12'd0942: exp <= 22'd3670333;
                12'd0943: exp <= 22'd3669269;
                12'd0944: exp <= 22'd3668204;
                12'd0945: exp <= 22'd3667138;
                12'd0946: exp <= 22'd3666071;
                12'd0947: exp <= 22'd3665003;
                12'd0948: exp <= 22'd3663935;
                12'd0949: exp <= 22'd3662865;
                12'd0950: exp <= 22'd3661794;
                12'd0951: exp <= 22'd3660723;
                12'd0952: exp <= 22'd3659650;
                12'd0953: exp <= 22'd3658577;
                12'd0954: exp <= 22'd3657503;
                12'd0955: exp <= 22'd3656428;
                12'd0956: exp <= 22'd3655352;
                12'd0957: exp <= 22'd3654275;
                12'd0958: exp <= 22'd3653197;
                12'd0959: exp <= 22'd3652118;
                12'd0960: exp <= 22'd3651038;
                12'd0961: exp <= 22'd3649957;
                12'd0962: exp <= 22'd3648876;
                12'd0963: exp <= 22'd3647793;
                12'd0964: exp <= 22'd3646710;
                12'd0965: exp <= 22'd3645626;
                12'd0966: exp <= 22'd3644541;
                12'd0967: exp <= 22'd3643454;
                12'd0968: exp <= 22'd3642367;
                12'd0969: exp <= 22'd3641279;
                12'd0970: exp <= 22'd3640191;
                12'd0971: exp <= 22'd3639101;
                12'd0972: exp <= 22'd3638010;
                12'd0973: exp <= 22'd3636919;
                12'd0974: exp <= 22'd3635826;
                12'd0975: exp <= 22'd3634733;
                12'd0976: exp <= 22'd3633638;
                12'd0977: exp <= 22'd3632543;
                12'd0978: exp <= 22'd3631447;
                12'd0979: exp <= 22'd3630350;
                12'd0980: exp <= 22'd3629252;
                12'd0981: exp <= 22'd3628153;
                12'd0982: exp <= 22'd3627054;
                12'd0983: exp <= 22'd3625953;
                12'd0984: exp <= 22'd3624852;
                12'd0985: exp <= 22'd3623749;
                12'd0986: exp <= 22'd3622646;
                12'd0987: exp <= 22'd3621542;
                12'd0988: exp <= 22'd3620437;
                12'd0989: exp <= 22'd3619331;
                12'd0990: exp <= 22'd3618224;
                12'd0991: exp <= 22'd3617116;
                12'd0992: exp <= 22'd3616007;
                12'd0993: exp <= 22'd3614898;
                12'd0994: exp <= 22'd3613787;
                12'd0995: exp <= 22'd3612676;
                12'd0996: exp <= 22'd3611564;
                12'd0997: exp <= 22'd3610450;
                12'd0998: exp <= 22'd3609336;
                12'd0999: exp <= 22'd3608222;
                12'd1000: exp <= 22'd3607106;
                12'd1001: exp <= 22'd3605989;
                12'd1002: exp <= 22'd3604871;
                12'd1003: exp <= 22'd3603753;
                12'd1004: exp <= 22'd3602634;
                12'd1005: exp <= 22'd3601513;
                12'd1006: exp <= 22'd3600392;
                12'd1007: exp <= 22'd3599270;
                12'd1008: exp <= 22'd3598147;
                12'd1009: exp <= 22'd3597024;
                12'd1010: exp <= 22'd3595899;
                12'd1011: exp <= 22'd3594773;
                12'd1012: exp <= 22'd3593647;
                12'd1013: exp <= 22'd3592520;
                12'd1014: exp <= 22'd3591391;
                12'd1015: exp <= 22'd3590262;
                12'd1016: exp <= 22'd3589132;
                12'd1017: exp <= 22'd3588002;
                12'd1018: exp <= 22'd3586870;
                12'd1019: exp <= 22'd3585737;
                12'd1020: exp <= 22'd3584604;
                12'd1021: exp <= 22'd3583470;
                12'd1022: exp <= 22'd3582334;
                12'd1023: exp <= 22'd3581198;
                12'd1024: exp <= 22'd3580061;
                12'd1025: exp <= 22'd3578924;
                12'd1026: exp <= 22'd3577785;
                12'd1027: exp <= 22'd3576645;
                12'd1028: exp <= 22'd3575505;
                12'd1029: exp <= 22'd3574364;
                12'd1030: exp <= 22'd3573221;
                12'd1031: exp <= 22'd3572078;
                12'd1032: exp <= 22'd3570935;
                12'd1033: exp <= 22'd3569790;
                12'd1034: exp <= 22'd3568644;
                12'd1035: exp <= 22'd3567498;
                12'd1036: exp <= 22'd3566350;
                12'd1037: exp <= 22'd3565202;
                12'd1038: exp <= 22'd3564053;
                12'd1039: exp <= 22'd3562903;
                12'd1040: exp <= 22'd3561752;
                12'd1041: exp <= 22'd3560600;
                12'd1042: exp <= 22'd3559448;
                12'd1043: exp <= 22'd3558295;
                12'd1044: exp <= 22'd3557140;
                12'd1045: exp <= 22'd3555985;
                12'd1046: exp <= 22'd3554829;
                12'd1047: exp <= 22'd3553672;
                12'd1048: exp <= 22'd3552515;
                12'd1049: exp <= 22'd3551356;
                12'd1050: exp <= 22'd3550197;
                12'd1051: exp <= 22'd3549036;
                12'd1052: exp <= 22'd3547875;
                12'd1053: exp <= 22'd3546713;
                12'd1054: exp <= 22'd3545551;
                12'd1055: exp <= 22'd3544387;
                12'd1056: exp <= 22'd3543222;
                12'd1057: exp <= 22'd3542057;
                12'd1058: exp <= 22'd3540891;
                12'd1059: exp <= 22'd3539724;
                12'd1060: exp <= 22'd3538556;
                12'd1061: exp <= 22'd3537387;
                12'd1062: exp <= 22'd3536217;
                12'd1063: exp <= 22'd3535047;
                12'd1064: exp <= 22'd3533876;
                12'd1065: exp <= 22'd3532703;
                12'd1066: exp <= 22'd3531530;
                12'd1067: exp <= 22'd3530357;
                12'd1068: exp <= 22'd3529182;
                12'd1069: exp <= 22'd3528006;
                12'd1070: exp <= 22'd3526830;
                12'd1071: exp <= 22'd3525653;
                12'd1072: exp <= 22'd3524475;
                12'd1073: exp <= 22'd3523296;
                12'd1074: exp <= 22'd3522116;
                12'd1075: exp <= 22'd3520936;
                12'd1076: exp <= 22'd3519754;
                12'd1077: exp <= 22'd3518572;
                12'd1078: exp <= 22'd3517389;
                12'd1079: exp <= 22'd3516205;
                12'd1080: exp <= 22'd3515020;
                12'd1081: exp <= 22'd3513835;
                12'd1082: exp <= 22'd3512648;
                12'd1083: exp <= 22'd3511461;
                12'd1084: exp <= 22'd3510273;
                12'd1085: exp <= 22'd3509084;
                12'd1086: exp <= 22'd3507894;
                12'd1087: exp <= 22'd3506704;
                12'd1088: exp <= 22'd3505512;
                12'd1089: exp <= 22'd3504320;
                12'd1090: exp <= 22'd3503127;
                12'd1091: exp <= 22'd3501933;
                12'd1092: exp <= 22'd3500738;
                12'd1093: exp <= 22'd3499543;
                12'd1094: exp <= 22'd3498346;
                12'd1095: exp <= 22'd3497149;
                12'd1096: exp <= 22'd3495951;
                12'd1097: exp <= 22'd3494752;
                12'd1098: exp <= 22'd3493553;
                12'd1099: exp <= 22'd3492352;
                12'd1100: exp <= 22'd3491151;
                12'd1101: exp <= 22'd3489949;
                12'd1102: exp <= 22'd3488746;
                12'd1103: exp <= 22'd3487542;
                12'd1104: exp <= 22'd3486338;
                12'd1105: exp <= 22'd3485132;
                12'd1106: exp <= 22'd3483926;
                12'd1107: exp <= 22'd3482719;
                12'd1108: exp <= 22'd3481511;
                12'd1109: exp <= 22'd3480302;
                12'd1110: exp <= 22'd3479093;
                12'd1111: exp <= 22'd3477883;
                12'd1112: exp <= 22'd3476672;
                12'd1113: exp <= 22'd3475460;
                12'd1114: exp <= 22'd3474247;
                12'd1115: exp <= 22'd3473033;
                12'd1116: exp <= 22'd3471819;
                12'd1117: exp <= 22'd3470604;
                12'd1118: exp <= 22'd3469388;
                12'd1119: exp <= 22'd3468171;
                12'd1120: exp <= 22'd3466954;
                12'd1121: exp <= 22'd3465735;
                12'd1122: exp <= 22'd3464516;
                12'd1123: exp <= 22'd3463296;
                12'd1124: exp <= 22'd3462075;
                12'd1125: exp <= 22'd3460854;
                12'd1126: exp <= 22'd3459631;
                12'd1127: exp <= 22'd3458408;
                12'd1128: exp <= 22'd3457184;
                12'd1129: exp <= 22'd3455959;
                12'd1130: exp <= 22'd3454734;
                12'd1131: exp <= 22'd3453508;
                12'd1132: exp <= 22'd3452280;
                12'd1133: exp <= 22'd3451052;
                12'd1134: exp <= 22'd3449824;
                12'd1135: exp <= 22'd3448594;
                12'd1136: exp <= 22'd3447364;
                12'd1137: exp <= 22'd3446132;
                12'd1138: exp <= 22'd3444900;
                12'd1139: exp <= 22'd3443668;
                12'd1140: exp <= 22'd3442434;
                12'd1141: exp <= 22'd3441200;
                12'd1142: exp <= 22'd3439965;
                12'd1143: exp <= 22'd3438729;
                12'd1144: exp <= 22'd3437492;
                12'd1145: exp <= 22'd3436255;
                12'd1146: exp <= 22'd3435016;
                12'd1147: exp <= 22'd3433777;
                12'd1148: exp <= 22'd3432537;
                12'd1149: exp <= 22'd3431297;
                12'd1150: exp <= 22'd3430055;
                12'd1151: exp <= 22'd3428813;
                12'd1152: exp <= 22'd3427570;
                12'd1153: exp <= 22'd3426326;
                12'd1154: exp <= 22'd3425082;
                12'd1155: exp <= 22'd3423836;
                12'd1156: exp <= 22'd3422590;
                12'd1157: exp <= 22'd3421343;
                12'd1158: exp <= 22'd3420096;
                12'd1159: exp <= 22'd3418847;
                12'd1160: exp <= 22'd3417598;
                12'd1161: exp <= 22'd3416348;
                12'd1162: exp <= 22'd3415097;
                12'd1163: exp <= 22'd3413846;
                12'd1164: exp <= 22'd3412593;
                12'd1165: exp <= 22'd3411340;
                12'd1166: exp <= 22'd3410086;
                12'd1167: exp <= 22'd3408832;
                12'd1168: exp <= 22'd3407576;
                12'd1169: exp <= 22'd3406320;
                12'd1170: exp <= 22'd3405063;
                12'd1171: exp <= 22'd3403805;
                12'd1172: exp <= 22'd3402547;
                12'd1173: exp <= 22'd3401288;
                12'd1174: exp <= 22'd3400028;
                12'd1175: exp <= 22'd3398767;
                12'd1176: exp <= 22'd3397505;
                12'd1177: exp <= 22'd3396243;
                12'd1178: exp <= 22'd3394980;
                12'd1179: exp <= 22'd3393716;
                12'd1180: exp <= 22'd3392451;
                12'd1181: exp <= 22'd3391186;
                12'd1182: exp <= 22'd3389920;
                12'd1183: exp <= 22'd3388653;
                12'd1184: exp <= 22'd3387385;
                12'd1185: exp <= 22'd3386117;
                12'd1186: exp <= 22'd3384848;
                12'd1187: exp <= 22'd3383578;
                12'd1188: exp <= 22'd3382307;
                12'd1189: exp <= 22'd3381035;
                12'd1190: exp <= 22'd3379763;
                12'd1191: exp <= 22'd3378490;
                12'd1192: exp <= 22'd3377217;
                12'd1193: exp <= 22'd3375942;
                12'd1194: exp <= 22'd3374667;
                12'd1195: exp <= 22'd3373391;
                12'd1196: exp <= 22'd3372114;
                12'd1197: exp <= 22'd3370837;
                12'd1198: exp <= 22'd3369558;
                12'd1199: exp <= 22'd3368279;
                12'd1200: exp <= 22'd3367000;
                12'd1201: exp <= 22'd3365719;
                12'd1202: exp <= 22'd3364438;
                12'd1203: exp <= 22'd3363156;
                12'd1204: exp <= 22'd3361873;
                12'd1205: exp <= 22'd3360590;
                12'd1206: exp <= 22'd3359306;
                12'd1207: exp <= 22'd3358021;
                12'd1208: exp <= 22'd3356735;
                12'd1209: exp <= 22'd3355449;
                12'd1210: exp <= 22'd3354161;
                12'd1211: exp <= 22'd3352874;
                12'd1212: exp <= 22'd3351585;
                12'd1213: exp <= 22'd3350296;
                12'd1214: exp <= 22'd3349005;
                12'd1215: exp <= 22'd3347715;
                12'd1216: exp <= 22'd3346423;
                12'd1217: exp <= 22'd3345131;
                12'd1218: exp <= 22'd3343838;
                12'd1219: exp <= 22'd3342544;
                12'd1220: exp <= 22'd3341249;
                12'd1221: exp <= 22'd3339954;
                12'd1222: exp <= 22'd3338658;
                12'd1223: exp <= 22'd3337361;
                12'd1224: exp <= 22'd3336064;
                12'd1225: exp <= 22'd3334766;
                12'd1226: exp <= 22'd3333467;
                12'd1227: exp <= 22'd3332167;
                12'd1228: exp <= 22'd3330867;
                12'd1229: exp <= 22'd3329566;
                12'd1230: exp <= 22'd3328264;
                12'd1231: exp <= 22'd3326961;
                12'd1232: exp <= 22'd3325658;
                12'd1233: exp <= 22'd3324354;
                12'd1234: exp <= 22'd3323049;
                12'd1235: exp <= 22'd3321744;
                12'd1236: exp <= 22'd3320438;
                12'd1237: exp <= 22'd3319131;
                12'd1238: exp <= 22'd3317823;
                12'd1239: exp <= 22'd3316515;
                12'd1240: exp <= 22'd3315206;
                12'd1241: exp <= 22'd3313896;
                12'd1242: exp <= 22'd3312586;
                12'd1243: exp <= 22'd3311275;
                12'd1244: exp <= 22'd3309963;
                12'd1245: exp <= 22'd3308650;
                12'd1246: exp <= 22'd3307337;
                12'd1247: exp <= 22'd3306023;
                12'd1248: exp <= 22'd3304708;
                12'd1249: exp <= 22'd3303393;
                12'd1250: exp <= 22'd3302077;
                12'd1251: exp <= 22'd3300760;
                12'd1252: exp <= 22'd3299442;
                12'd1253: exp <= 22'd3298124;
                12'd1254: exp <= 22'd3296805;
                12'd1255: exp <= 22'd3295485;
                12'd1256: exp <= 22'd3294165;
                12'd1257: exp <= 22'd3292844;
                12'd1258: exp <= 22'd3291522;
                12'd1259: exp <= 22'd3290200;
                12'd1260: exp <= 22'd3288876;
                12'd1261: exp <= 22'd3287552;
                12'd1262: exp <= 22'd3286228;
                12'd1263: exp <= 22'd3284903;
                12'd1264: exp <= 22'd3283577;
                12'd1265: exp <= 22'd3282250;
                12'd1266: exp <= 22'd3280923;
                12'd1267: exp <= 22'd3279594;
                12'd1268: exp <= 22'd3278266;
                12'd1269: exp <= 22'd3276936;
                12'd1270: exp <= 22'd3275606;
                12'd1271: exp <= 22'd3274275;
                12'd1272: exp <= 22'd3272944;
                12'd1273: exp <= 22'd3271611;
                12'd1274: exp <= 22'd3270278;
                12'd1275: exp <= 22'd3268945;
                12'd1276: exp <= 22'd3267610;
                12'd1277: exp <= 22'd3266275;
                12'd1278: exp <= 22'd3264940;
                12'd1279: exp <= 22'd3263603;
                12'd1280: exp <= 22'd3262266;
                12'd1281: exp <= 22'd3260928;
                12'd1282: exp <= 22'd3259590;
                12'd1283: exp <= 22'd3258251;
                12'd1284: exp <= 22'd3256911;
                12'd1285: exp <= 22'd3255571;
                12'd1286: exp <= 22'd3254229;
                12'd1287: exp <= 22'd3252888;
                12'd1288: exp <= 22'd3251545;
                12'd1289: exp <= 22'd3250202;
                12'd1290: exp <= 22'd3248858;
                12'd1291: exp <= 22'd3247513;
                12'd1292: exp <= 22'd3246168;
                12'd1293: exp <= 22'd3244822;
                12'd1294: exp <= 22'd3243476;
                12'd1295: exp <= 22'd3242128;
                12'd1296: exp <= 22'd3240780;
                12'd1297: exp <= 22'd3239432;
                12'd1298: exp <= 22'd3238082;
                12'd1299: exp <= 22'd3236733;
                12'd1300: exp <= 22'd3235382;
                12'd1301: exp <= 22'd3234031;
                12'd1302: exp <= 22'd3232679;
                12'd1303: exp <= 22'd3231326;
                12'd1304: exp <= 22'd3229973;
                12'd1305: exp <= 22'd3228619;
                12'd1306: exp <= 22'd3227264;
                12'd1307: exp <= 22'd3225909;
                12'd1308: exp <= 22'd3224553;
                12'd1309: exp <= 22'd3223196;
                12'd1310: exp <= 22'd3221839;
                12'd1311: exp <= 22'd3220481;
                12'd1312: exp <= 22'd3219122;
                12'd1313: exp <= 22'd3217763;
                12'd1314: exp <= 22'd3216403;
                12'd1315: exp <= 22'd3215043;
                12'd1316: exp <= 22'd3213681;
                12'd1317: exp <= 22'd3212319;
                12'd1318: exp <= 22'd3210957;
                12'd1319: exp <= 22'd3209594;
                12'd1320: exp <= 22'd3208230;
                12'd1321: exp <= 22'd3206865;
                12'd1322: exp <= 22'd3205500;
                12'd1323: exp <= 22'd3204134;
                12'd1324: exp <= 22'd3202768;
                12'd1325: exp <= 22'd3201401;
                12'd1326: exp <= 22'd3200033;
                12'd1327: exp <= 22'd3198664;
                12'd1328: exp <= 22'd3197295;
                12'd1329: exp <= 22'd3195926;
                12'd1330: exp <= 22'd3194555;
                12'd1331: exp <= 22'd3193184;
                12'd1332: exp <= 22'd3191813;
                12'd1333: exp <= 22'd3190440;
                12'd1334: exp <= 22'd3189067;
                12'd1335: exp <= 22'd3187694;
                12'd1336: exp <= 22'd3186319;
                12'd1337: exp <= 22'd3184945;
                12'd1338: exp <= 22'd3183569;
                12'd1339: exp <= 22'd3182193;
                12'd1340: exp <= 22'd3180816;
                12'd1341: exp <= 22'd3179439;
                12'd1342: exp <= 22'd3178061;
                12'd1343: exp <= 22'd3176682;
                12'd1344: exp <= 22'd3175303;
                12'd1345: exp <= 22'd3173923;
                12'd1346: exp <= 22'd3172542;
                12'd1347: exp <= 22'd3171161;
                12'd1348: exp <= 22'd3169779;
                12'd1349: exp <= 22'd3168396;
                12'd1350: exp <= 22'd3167013;
                12'd1351: exp <= 22'd3165630;
                12'd1352: exp <= 22'd3164245;
                12'd1353: exp <= 22'd3162860;
                12'd1354: exp <= 22'd3161474;
                12'd1355: exp <= 22'd3160088;
                12'd1356: exp <= 22'd3158701;
                12'd1357: exp <= 22'd3157314;
                12'd1358: exp <= 22'd3155926;
                12'd1359: exp <= 22'd3154537;
                12'd1360: exp <= 22'd3153148;
                12'd1361: exp <= 22'd3151758;
                12'd1362: exp <= 22'd3150367;
                12'd1363: exp <= 22'd3148976;
                12'd1364: exp <= 22'd3147584;
                12'd1365: exp <= 22'd3146191;
                12'd1366: exp <= 22'd3144798;
                12'd1367: exp <= 22'd3143404;
                12'd1368: exp <= 22'd3142010;
                12'd1369: exp <= 22'd3140615;
                12'd1370: exp <= 22'd3139220;
                12'd1371: exp <= 22'd3137823;
                12'd1372: exp <= 22'd3136427;
                12'd1373: exp <= 22'd3135029;
                12'd1374: exp <= 22'd3133631;
                12'd1375: exp <= 22'd3132233;
                12'd1376: exp <= 22'd3130833;
                12'd1377: exp <= 22'd3129434;
                12'd1378: exp <= 22'd3128033;
                12'd1379: exp <= 22'd3126632;
                12'd1380: exp <= 22'd3125230;
                12'd1381: exp <= 22'd3123828;
                12'd1382: exp <= 22'd3122425;
                12'd1383: exp <= 22'd3121022;
                12'd1384: exp <= 22'd3119618;
                12'd1385: exp <= 22'd3118213;
                12'd1386: exp <= 22'd3116808;
                12'd1387: exp <= 22'd3115402;
                12'd1388: exp <= 22'd3113996;
                12'd1389: exp <= 22'd3112588;
                12'd1390: exp <= 22'd3111181;
                12'd1391: exp <= 22'd3109773;
                12'd1392: exp <= 22'd3108364;
                12'd1393: exp <= 22'd3106954;
                12'd1394: exp <= 22'd3105544;
                12'd1395: exp <= 22'd3104134;
                12'd1396: exp <= 22'd3102722;
                12'd1397: exp <= 22'd3101310;
                12'd1398: exp <= 22'd3099898;
                12'd1399: exp <= 22'd3098485;
                12'd1400: exp <= 22'd3097071;
                12'd1401: exp <= 22'd3095657;
                12'd1402: exp <= 22'd3094243;
                12'd1403: exp <= 22'd3092827;
                12'd1404: exp <= 22'd3091411;
                12'd1405: exp <= 22'd3089995;
                12'd1406: exp <= 22'd3088578;
                12'd1407: exp <= 22'd3087160;
                12'd1408: exp <= 22'd3085742;
                12'd1409: exp <= 22'd3084323;
                12'd1410: exp <= 22'd3082903;
                12'd1411: exp <= 22'd3081483;
                12'd1412: exp <= 22'd3080063;
                12'd1413: exp <= 22'd3078642;
                12'd1414: exp <= 22'd3077220;
                12'd1415: exp <= 22'd3075797;
                12'd1416: exp <= 22'd3074375;
                12'd1417: exp <= 22'd3072951;
                12'd1418: exp <= 22'd3071527;
                12'd1419: exp <= 22'd3070102;
                12'd1420: exp <= 22'd3068677;
                12'd1421: exp <= 22'd3067251;
                12'd1422: exp <= 22'd3065825;
                12'd1423: exp <= 22'd3064398;
                12'd1424: exp <= 22'd3062971;
                12'd1425: exp <= 22'd3061543;
                12'd1426: exp <= 22'd3060114;
                12'd1427: exp <= 22'd3058685;
                12'd1428: exp <= 22'd3057255;
                12'd1429: exp <= 22'd3055825;
                12'd1430: exp <= 22'd3054394;
                12'd1431: exp <= 22'd3052962;
                12'd1432: exp <= 22'd3051530;
                12'd1433: exp <= 22'd3050098;
                12'd1434: exp <= 22'd3048665;
                12'd1435: exp <= 22'd3047231;
                12'd1436: exp <= 22'd3045797;
                12'd1437: exp <= 22'd3044362;
                12'd1438: exp <= 22'd3042927;
                12'd1439: exp <= 22'd3041491;
                12'd1440: exp <= 22'd3040054;
                12'd1441: exp <= 22'd3038617;
                12'd1442: exp <= 22'd3037180;
                12'd1443: exp <= 22'd3035742;
                12'd1444: exp <= 22'd3034303;
                12'd1445: exp <= 22'd3032864;
                12'd1446: exp <= 22'd3031424;
                12'd1447: exp <= 22'd3029984;
                12'd1448: exp <= 22'd3028543;
                12'd1449: exp <= 22'd3027101;
                12'd1450: exp <= 22'd3025659;
                12'd1451: exp <= 22'd3024217;
                12'd1452: exp <= 22'd3022774;
                12'd1453: exp <= 22'd3021330;
                12'd1454: exp <= 22'd3019886;
                12'd1455: exp <= 22'd3018441;
                12'd1456: exp <= 22'd3016996;
                12'd1457: exp <= 22'd3015550;
                12'd1458: exp <= 22'd3014104;
                12'd1459: exp <= 22'd3012657;
                12'd1460: exp <= 22'd3011210;
                12'd1461: exp <= 22'd3009762;
                12'd1462: exp <= 22'd3008313;
                12'd1463: exp <= 22'd3006864;
                12'd1464: exp <= 22'd3005415;
                12'd1465: exp <= 22'd3003964;
                12'd1466: exp <= 22'd3002514;
                12'd1467: exp <= 22'd3001063;
                12'd1468: exp <= 22'd2999611;
                12'd1469: exp <= 22'd2998159;
                12'd1470: exp <= 22'd2996706;
                12'd1471: exp <= 22'd2995253;
                12'd1472: exp <= 22'd2993799;
                12'd1473: exp <= 22'd2992345;
                12'd1474: exp <= 22'd2990890;
                12'd1475: exp <= 22'd2989434;
                12'd1476: exp <= 22'd2987979;
                12'd1477: exp <= 22'd2986522;
                12'd1478: exp <= 22'd2985065;
                12'd1479: exp <= 22'd2983608;
                12'd1480: exp <= 22'd2982150;
                12'd1481: exp <= 22'd2980691;
                12'd1482: exp <= 22'd2979232;
                12'd1483: exp <= 22'd2977773;
                12'd1484: exp <= 22'd2976313;
                12'd1485: exp <= 22'd2974852;
                12'd1486: exp <= 22'd2973391;
                12'd1487: exp <= 22'd2971929;
                12'd1488: exp <= 22'd2970467;
                12'd1489: exp <= 22'd2969004;
                12'd1490: exp <= 22'd2967541;
                12'd1491: exp <= 22'd2966078;
                12'd1492: exp <= 22'd2964613;
                12'd1493: exp <= 22'd2963149;
                12'd1494: exp <= 22'd2961684;
                12'd1495: exp <= 22'd2960218;
                12'd1496: exp <= 22'd2958752;
                12'd1497: exp <= 22'd2957285;
                12'd1498: exp <= 22'd2955818;
                12'd1499: exp <= 22'd2954350;
                12'd1500: exp <= 22'd2952882;
                12'd1501: exp <= 22'd2951413;
                12'd1502: exp <= 22'd2949944;
                12'd1503: exp <= 22'd2948474;
                12'd1504: exp <= 22'd2947004;
                12'd1505: exp <= 22'd2945533;
                12'd1506: exp <= 22'd2944062;
                12'd1507: exp <= 22'd2942590;
                12'd1508: exp <= 22'd2941118;
                12'd1509: exp <= 22'd2939645;
                12'd1510: exp <= 22'd2938172;
                12'd1511: exp <= 22'd2936698;
                12'd1512: exp <= 22'd2935224;
                12'd1513: exp <= 22'd2933749;
                12'd1514: exp <= 22'd2932274;
                12'd1515: exp <= 22'd2930798;
                12'd1516: exp <= 22'd2929322;
                12'd1517: exp <= 22'd2927845;
                12'd1518: exp <= 22'd2926368;
                12'd1519: exp <= 22'd2924890;
                12'd1520: exp <= 22'd2923412;
                12'd1521: exp <= 22'd2921934;
                12'd1522: exp <= 22'd2920454;
                12'd1523: exp <= 22'd2918975;
                12'd1524: exp <= 22'd2917495;
                12'd1525: exp <= 22'd2916014;
                12'd1526: exp <= 22'd2914533;
                12'd1527: exp <= 22'd2913052;
                12'd1528: exp <= 22'd2911570;
                12'd1529: exp <= 22'd2910087;
                12'd1530: exp <= 22'd2908604;
                12'd1531: exp <= 22'd2907121;
                12'd1532: exp <= 22'd2905637;
                12'd1533: exp <= 22'd2904152;
                12'd1534: exp <= 22'd2902667;
                12'd1535: exp <= 22'd2901182;
                12'd1536: exp <= 22'd2899696;
                12'd1537: exp <= 22'd2898210;
                12'd1538: exp <= 22'd2896723;
                12'd1539: exp <= 22'd2895236;
                12'd1540: exp <= 22'd2893748;
                12'd1541: exp <= 22'd2892260;
                12'd1542: exp <= 22'd2890772;
                12'd1543: exp <= 22'd2889282;
                12'd1544: exp <= 22'd2887793;
                12'd1545: exp <= 22'd2886303;
                12'd1546: exp <= 22'd2884812;
                12'd1547: exp <= 22'd2883321;
                12'd1548: exp <= 22'd2881830;
                12'd1549: exp <= 22'd2880338;
                12'd1550: exp <= 22'd2878846;
                12'd1551: exp <= 22'd2877353;
                12'd1552: exp <= 22'd2875860;
                12'd1553: exp <= 22'd2874366;
                12'd1554: exp <= 22'd2872872;
                12'd1555: exp <= 22'd2871377;
                12'd1556: exp <= 22'd2869882;
                12'd1557: exp <= 22'd2868386;
                12'd1558: exp <= 22'd2866890;
                12'd1559: exp <= 22'd2865394;
                12'd1560: exp <= 22'd2863897;
                12'd1561: exp <= 22'd2862400;
                12'd1562: exp <= 22'd2860902;
                12'd1563: exp <= 22'd2859404;
                12'd1564: exp <= 22'd2857905;
                12'd1565: exp <= 22'd2856406;
                12'd1566: exp <= 22'd2854906;
                12'd1567: exp <= 22'd2853406;
                12'd1568: exp <= 22'd2851906;
                12'd1569: exp <= 22'd2850405;
                12'd1570: exp <= 22'd2848903;
                12'd1571: exp <= 22'd2847401;
                12'd1572: exp <= 22'd2845899;
                12'd1573: exp <= 22'd2844396;
                12'd1574: exp <= 22'd2842893;
                12'd1575: exp <= 22'd2841390;
                12'd1576: exp <= 22'd2839886;
                12'd1577: exp <= 22'd2838381;
                12'd1578: exp <= 22'd2836876;
                12'd1579: exp <= 22'd2835371;
                12'd1580: exp <= 22'd2833865;
                12'd1581: exp <= 22'd2832359;
                12'd1582: exp <= 22'd2830852;
                12'd1583: exp <= 22'd2829345;
                12'd1584: exp <= 22'd2827838;
                12'd1585: exp <= 22'd2826330;
                12'd1586: exp <= 22'd2824822;
                12'd1587: exp <= 22'd2823313;
                12'd1588: exp <= 22'd2821804;
                12'd1589: exp <= 22'd2820294;
                12'd1590: exp <= 22'd2818784;
                12'd1591: exp <= 22'd2817274;
                12'd1592: exp <= 22'd2815763;
                12'd1593: exp <= 22'd2814251;
                12'd1594: exp <= 22'd2812740;
                12'd1595: exp <= 22'd2811227;
                12'd1596: exp <= 22'd2809715;
                12'd1597: exp <= 22'd2808202;
                12'd1598: exp <= 22'd2806688;
                12'd1599: exp <= 22'd2805174;
                12'd1600: exp <= 22'd2803660;
                12'd1601: exp <= 22'd2802146;
                12'd1602: exp <= 22'd2800630;
                12'd1603: exp <= 22'd2799115;
                12'd1604: exp <= 22'd2797599;
                12'd1605: exp <= 22'd2796083;
                12'd1606: exp <= 22'd2794566;
                12'd1607: exp <= 22'd2793049;
                12'd1608: exp <= 22'd2791531;
                12'd1609: exp <= 22'd2790013;
                12'd1610: exp <= 22'd2788495;
                12'd1611: exp <= 22'd2786976;
                12'd1612: exp <= 22'd2785457;
                12'd1613: exp <= 22'd2783937;
                12'd1614: exp <= 22'd2782417;
                12'd1615: exp <= 22'd2780897;
                12'd1616: exp <= 22'd2779376;
                12'd1617: exp <= 22'd2777855;
                12'd1618: exp <= 22'd2776333;
                12'd1619: exp <= 22'd2774811;
                12'd1620: exp <= 22'd2773289;
                12'd1621: exp <= 22'd2771766;
                12'd1622: exp <= 22'd2770243;
                12'd1623: exp <= 22'd2768719;
                12'd1624: exp <= 22'd2767195;
                12'd1625: exp <= 22'd2765671;
                12'd1626: exp <= 22'd2764146;
                12'd1627: exp <= 22'd2762621;
                12'd1628: exp <= 22'd2761095;
                12'd1629: exp <= 22'd2759569;
                12'd1630: exp <= 22'd2758043;
                12'd1631: exp <= 22'd2756516;
                12'd1632: exp <= 22'd2754989;
                12'd1633: exp <= 22'd2753462;
                12'd1634: exp <= 22'd2751934;
                12'd1635: exp <= 22'd2750406;
                12'd1636: exp <= 22'd2748877;
                12'd1637: exp <= 22'd2747348;
                12'd1638: exp <= 22'd2745818;
                12'd1639: exp <= 22'd2744289;
                12'd1640: exp <= 22'd2742758;
                12'd1641: exp <= 22'd2741228;
                12'd1642: exp <= 22'd2739697;
                12'd1643: exp <= 22'd2738166;
                12'd1644: exp <= 22'd2736634;
                12'd1645: exp <= 22'd2735102;
                12'd1646: exp <= 22'd2733569;
                12'd1647: exp <= 22'd2732037;
                12'd1648: exp <= 22'd2730503;
                12'd1649: exp <= 22'd2728970;
                12'd1650: exp <= 22'd2727436;
                12'd1651: exp <= 22'd2725902;
                12'd1652: exp <= 22'd2724367;
                12'd1653: exp <= 22'd2722832;
                12'd1654: exp <= 22'd2721296;
                12'd1655: exp <= 22'd2719761;
                12'd1656: exp <= 22'd2718224;
                12'd1657: exp <= 22'd2716688;
                12'd1658: exp <= 22'd2715151;
                12'd1659: exp <= 22'd2713614;
                12'd1660: exp <= 22'd2712076;
                12'd1661: exp <= 22'd2710538;
                12'd1662: exp <= 22'd2709000;
                12'd1663: exp <= 22'd2707461;
                12'd1664: exp <= 22'd2705922;
                12'd1665: exp <= 22'd2704383;
                12'd1666: exp <= 22'd2702843;
                12'd1667: exp <= 22'd2701303;
                12'd1668: exp <= 22'd2699762;
                12'd1669: exp <= 22'd2698221;
                12'd1670: exp <= 22'd2696680;
                12'd1671: exp <= 22'd2695139;
                12'd1672: exp <= 22'd2693597;
                12'd1673: exp <= 22'd2692055;
                12'd1674: exp <= 22'd2690512;
                12'd1675: exp <= 22'd2688969;
                12'd1676: exp <= 22'd2687426;
                12'd1677: exp <= 22'd2685882;
                12'd1678: exp <= 22'd2684338;
                12'd1679: exp <= 22'd2682794;
                12'd1680: exp <= 22'd2681249;
                12'd1681: exp <= 22'd2679704;
                12'd1682: exp <= 22'd2678159;
                12'd1683: exp <= 22'd2676613;
                12'd1684: exp <= 22'd2675067;
                12'd1685: exp <= 22'd2673521;
                12'd1686: exp <= 22'd2671974;
                12'd1687: exp <= 22'd2670427;
                12'd1688: exp <= 22'd2668879;
                12'd1689: exp <= 22'd2667332;
                12'd1690: exp <= 22'd2665784;
                12'd1691: exp <= 22'd2664235;
                12'd1692: exp <= 22'd2662686;
                12'd1693: exp <= 22'd2661137;
                12'd1694: exp <= 22'd2659588;
                12'd1695: exp <= 22'd2658038;
                12'd1696: exp <= 22'd2656488;
                12'd1697: exp <= 22'd2654938;
                12'd1698: exp <= 22'd2653387;
                12'd1699: exp <= 22'd2651836;
                12'd1700: exp <= 22'd2650285;
                12'd1701: exp <= 22'd2648733;
                12'd1702: exp <= 22'd2647181;
                12'd1703: exp <= 22'd2645629;
                12'd1704: exp <= 22'd2644076;
                12'd1705: exp <= 22'd2642523;
                12'd1706: exp <= 22'd2640970;
                12'd1707: exp <= 22'd2639416;
                12'd1708: exp <= 22'd2637862;
                12'd1709: exp <= 22'd2636308;
                12'd1710: exp <= 22'd2634753;
                12'd1711: exp <= 22'd2633198;
                12'd1712: exp <= 22'd2631643;
                12'd1713: exp <= 22'd2630087;
                12'd1714: exp <= 22'd2628532;
                12'd1715: exp <= 22'd2626975;
                12'd1716: exp <= 22'd2625419;
                12'd1717: exp <= 22'd2623862;
                12'd1718: exp <= 22'd2622305;
                12'd1719: exp <= 22'd2620748;
                12'd1720: exp <= 22'd2619190;
                12'd1721: exp <= 22'd2617632;
                12'd1722: exp <= 22'd2616074;
                12'd1723: exp <= 22'd2614515;
                12'd1724: exp <= 22'd2612956;
                12'd1725: exp <= 22'd2611397;
                12'd1726: exp <= 22'd2609837;
                12'd1727: exp <= 22'd2608278;
                12'd1728: exp <= 22'd2606717;
                12'd1729: exp <= 22'd2605157;
                12'd1730: exp <= 22'd2603596;
                12'd1731: exp <= 22'd2602035;
                12'd1732: exp <= 22'd2600474;
                12'd1733: exp <= 22'd2598912;
                12'd1734: exp <= 22'd2597350;
                12'd1735: exp <= 22'd2595788;
                12'd1736: exp <= 22'd2594226;
                12'd1737: exp <= 22'd2592663;
                12'd1738: exp <= 22'd2591100;
                12'd1739: exp <= 22'd2589536;
                12'd1740: exp <= 22'd2587973;
                12'd1741: exp <= 22'd2586409;
                12'd1742: exp <= 22'd2584844;
                12'd1743: exp <= 22'd2583280;
                12'd1744: exp <= 22'd2581715;
                12'd1745: exp <= 22'd2580150;
                12'd1746: exp <= 22'd2578584;
                12'd1747: exp <= 22'd2577019;
                12'd1748: exp <= 22'd2575453;
                12'd1749: exp <= 22'd2573887;
                12'd1750: exp <= 22'd2572320;
                12'd1751: exp <= 22'd2570753;
                12'd1752: exp <= 22'd2569186;
                12'd1753: exp <= 22'd2567619;
                12'd1754: exp <= 22'd2566051;
                12'd1755: exp <= 22'd2564483;
                12'd1756: exp <= 22'd2562915;
                12'd1757: exp <= 22'd2561347;
                12'd1758: exp <= 22'd2559778;
                12'd1759: exp <= 22'd2558209;
                12'd1760: exp <= 22'd2556640;
                12'd1761: exp <= 22'd2555070;
                12'd1762: exp <= 22'd2553500;
                12'd1763: exp <= 22'd2551930;
                12'd1764: exp <= 22'd2550360;
                12'd1765: exp <= 22'd2548789;
                12'd1766: exp <= 22'd2547218;
                12'd1767: exp <= 22'd2545647;
                12'd1768: exp <= 22'd2544076;
                12'd1769: exp <= 22'd2542504;
                12'd1770: exp <= 22'd2540932;
                12'd1771: exp <= 22'd2539360;
                12'd1772: exp <= 22'd2537787;
                12'd1773: exp <= 22'd2536215;
                12'd1774: exp <= 22'd2534642;
                12'd1775: exp <= 22'd2533069;
                12'd1776: exp <= 22'd2531495;
                12'd1777: exp <= 22'd2529921;
                12'd1778: exp <= 22'd2528347;
                12'd1779: exp <= 22'd2526773;
                12'd1780: exp <= 22'd2525199;
                12'd1781: exp <= 22'd2523624;
                12'd1782: exp <= 22'd2522049;
                12'd1783: exp <= 22'd2520473;
                12'd1784: exp <= 22'd2518898;
                12'd1785: exp <= 22'd2517322;
                12'd1786: exp <= 22'd2515746;
                12'd1787: exp <= 22'd2514170;
                12'd1788: exp <= 22'd2512593;
                12'd1789: exp <= 22'd2511017;
                12'd1790: exp <= 22'd2509440;
                12'd1791: exp <= 22'd2507863;
                12'd1792: exp <= 22'd2506285;
                12'd1793: exp <= 22'd2504707;
                12'd1794: exp <= 22'd2503129;
                12'd1795: exp <= 22'd2501551;
                12'd1796: exp <= 22'd2499973;
                12'd1797: exp <= 22'd2498394;
                12'd1798: exp <= 22'd2496815;
                12'd1799: exp <= 22'd2495236;
                12'd1800: exp <= 22'd2493657;
                12'd1801: exp <= 22'd2492077;
                12'd1802: exp <= 22'd2490497;
                12'd1803: exp <= 22'd2488917;
                12'd1804: exp <= 22'd2487337;
                12'd1805: exp <= 22'd2485756;
                12'd1806: exp <= 22'd2484176;
                12'd1807: exp <= 22'd2482595;
                12'd1808: exp <= 22'd2481013;
                12'd1809: exp <= 22'd2479432;
                12'd1810: exp <= 22'd2477850;
                12'd1811: exp <= 22'd2476268;
                12'd1812: exp <= 22'd2474686;
                12'd1813: exp <= 22'd2473104;
                12'd1814: exp <= 22'd2471522;
                12'd1815: exp <= 22'd2469939;
                12'd1816: exp <= 22'd2468356;
                12'd1817: exp <= 22'd2466773;
                12'd1818: exp <= 22'd2465189;
                12'd1819: exp <= 22'd2463605;
                12'd1820: exp <= 22'd2462022;
                12'd1821: exp <= 22'd2460438;
                12'd1822: exp <= 22'd2458853;
                12'd1823: exp <= 22'd2457269;
                12'd1824: exp <= 22'd2455684;
                12'd1825: exp <= 22'd2454099;
                12'd1826: exp <= 22'd2452514;
                12'd1827: exp <= 22'd2450929;
                12'd1828: exp <= 22'd2449343;
                12'd1829: exp <= 22'd2447757;
                12'd1830: exp <= 22'd2446171;
                12'd1831: exp <= 22'd2444585;
                12'd1832: exp <= 22'd2442999;
                12'd1833: exp <= 22'd2441412;
                12'd1834: exp <= 22'd2439826;
                12'd1835: exp <= 22'd2438239;
                12'd1836: exp <= 22'd2436651;
                12'd1837: exp <= 22'd2435064;
                12'd1838: exp <= 22'd2433476;
                12'd1839: exp <= 22'd2431889;
                12'd1840: exp <= 22'd2430301;
                12'd1841: exp <= 22'd2428713;
                12'd1842: exp <= 22'd2427124;
                12'd1843: exp <= 22'd2425536;
                12'd1844: exp <= 22'd2423947;
                12'd1845: exp <= 22'd2422358;
                12'd1846: exp <= 22'd2420769;
                12'd1847: exp <= 22'd2419179;
                12'd1848: exp <= 22'd2417590;
                12'd1849: exp <= 22'd2416000;
                12'd1850: exp <= 22'd2414410;
                12'd1851: exp <= 22'd2412820;
                12'd1852: exp <= 22'd2411230;
                12'd1853: exp <= 22'd2409640;
                12'd1854: exp <= 22'd2408049;
                12'd1855: exp <= 22'd2406458;
                12'd1856: exp <= 22'd2404867;
                12'd1857: exp <= 22'd2403276;
                12'd1858: exp <= 22'd2401685;
                12'd1859: exp <= 22'd2400093;
                12'd1860: exp <= 22'd2398501;
                12'd1861: exp <= 22'd2396909;
                12'd1862: exp <= 22'd2395317;
                12'd1863: exp <= 22'd2393725;
                12'd1864: exp <= 22'd2392133;
                12'd1865: exp <= 22'd2390540;
                12'd1866: exp <= 22'd2388947;
                12'd1867: exp <= 22'd2387354;
                12'd1868: exp <= 22'd2385761;
                12'd1869: exp <= 22'd2384168;
                12'd1870: exp <= 22'd2382575;
                12'd1871: exp <= 22'd2380981;
                12'd1872: exp <= 22'd2379387;
                12'd1873: exp <= 22'd2377793;
                12'd1874: exp <= 22'd2376199;
                12'd1875: exp <= 22'd2374605;
                12'd1876: exp <= 22'd2373010;
                12'd1877: exp <= 22'd2371416;
                12'd1878: exp <= 22'd2369821;
                12'd1879: exp <= 22'd2368226;
                12'd1880: exp <= 22'd2366631;
                12'd1881: exp <= 22'd2365036;
                12'd1882: exp <= 22'd2363440;
                12'd1883: exp <= 22'd2361845;
                12'd1884: exp <= 22'd2360249;
                12'd1885: exp <= 22'd2358653;
                12'd1886: exp <= 22'd2357057;
                12'd1887: exp <= 22'd2355461;
                12'd1888: exp <= 22'd2353865;
                12'd1889: exp <= 22'd2352268;
                12'd1890: exp <= 22'd2350672;
                12'd1891: exp <= 22'd2349075;
                12'd1892: exp <= 22'd2347478;
                12'd1893: exp <= 22'd2345881;
                12'd1894: exp <= 22'd2344284;
                12'd1895: exp <= 22'd2342686;
                12'd1896: exp <= 22'd2341089;
                12'd1897: exp <= 22'd2339491;
                12'd1898: exp <= 22'd2337893;
                12'd1899: exp <= 22'd2336295;
                12'd1900: exp <= 22'd2334697;
                12'd1901: exp <= 22'd2333099;
                12'd1902: exp <= 22'd2331501;
                12'd1903: exp <= 22'd2329902;
                12'd1904: exp <= 22'd2328304;
                12'd1905: exp <= 22'd2326705;
                12'd1906: exp <= 22'd2325106;
                12'd1907: exp <= 22'd2323507;
                12'd1908: exp <= 22'd2321908;
                12'd1909: exp <= 22'd2320309;
                12'd1910: exp <= 22'd2318709;
                12'd1911: exp <= 22'd2317110;
                12'd1912: exp <= 22'd2315510;
                12'd1913: exp <= 22'd2313910;
                12'd1914: exp <= 22'd2312310;
                12'd1915: exp <= 22'd2310710;
                12'd1916: exp <= 22'd2309110;
                12'd1917: exp <= 22'd2307510;
                12'd1918: exp <= 22'd2305909;
                12'd1919: exp <= 22'd2304309;
                12'd1920: exp <= 22'd2302708;
                12'd1921: exp <= 22'd2301107;
                12'd1922: exp <= 22'd2299506;
                12'd1923: exp <= 22'd2297905;
                12'd1924: exp <= 22'd2296304;
                12'd1925: exp <= 22'd2294703;
                12'd1926: exp <= 22'd2293101;
                12'd1927: exp <= 22'd2291500;
                12'd1928: exp <= 22'd2289898;
                12'd1929: exp <= 22'd2288296;
                12'd1930: exp <= 22'd2286694;
                12'd1931: exp <= 22'd2285092;
                12'd1932: exp <= 22'd2283490;
                12'd1933: exp <= 22'd2281888;
                12'd1934: exp <= 22'd2280286;
                12'd1935: exp <= 22'd2278684;
                12'd1936: exp <= 22'd2277081;
                12'd1937: exp <= 22'd2275478;
                12'd1938: exp <= 22'd2273876;
                12'd1939: exp <= 22'd2272273;
                12'd1940: exp <= 22'd2270670;
                12'd1941: exp <= 22'd2269067;
                12'd1942: exp <= 22'd2267464;
                12'd1943: exp <= 22'd2265861;
                12'd1944: exp <= 22'd2264257;
                12'd1945: exp <= 22'd2262654;
                12'd1946: exp <= 22'd2261050;
                12'd1947: exp <= 22'd2259447;
                12'd1948: exp <= 22'd2257843;
                12'd1949: exp <= 22'd2256239;
                12'd1950: exp <= 22'd2254635;
                12'd1951: exp <= 22'd2253031;
                12'd1952: exp <= 22'd2251427;
                12'd1953: exp <= 22'd2249823;
                12'd1954: exp <= 22'd2248219;
                12'd1955: exp <= 22'd2246614;
                12'd1956: exp <= 22'd2245010;
                12'd1957: exp <= 22'd2243405;
                12'd1958: exp <= 22'd2241801;
                12'd1959: exp <= 22'd2240196;
                12'd1960: exp <= 22'd2238591;
                12'd1961: exp <= 22'd2236986;
                12'd1962: exp <= 22'd2235381;
                12'd1963: exp <= 22'd2233776;
                12'd1964: exp <= 22'd2232171;
                12'd1965: exp <= 22'd2230566;
                12'd1966: exp <= 22'd2228961;
                12'd1967: exp <= 22'd2227355;
                12'd1968: exp <= 22'd2225750;
                12'd1969: exp <= 22'd2224144;
                12'd1970: exp <= 22'd2222539;
                12'd1971: exp <= 22'd2220933;
                12'd1972: exp <= 22'd2219327;
                12'd1973: exp <= 22'd2217722;
                12'd1974: exp <= 22'd2216116;
                12'd1975: exp <= 22'd2214510;
                12'd1976: exp <= 22'd2212904;
                12'd1977: exp <= 22'd2211298;
                12'd1978: exp <= 22'd2209692;
                12'd1979: exp <= 22'd2208085;
                12'd1980: exp <= 22'd2206479;
                12'd1981: exp <= 22'd2204873;
                12'd1982: exp <= 22'd2203266;
                12'd1983: exp <= 22'd2201660;
                12'd1984: exp <= 22'd2200053;
                12'd1985: exp <= 22'd2198447;
                12'd1986: exp <= 22'd2196840;
                12'd1987: exp <= 22'd2195233;
                12'd1988: exp <= 22'd2193627;
                12'd1989: exp <= 22'd2192020;
                12'd1990: exp <= 22'd2190413;
                12'd1991: exp <= 22'd2188806;
                12'd1992: exp <= 22'd2187199;
                12'd1993: exp <= 22'd2185592;
                12'd1994: exp <= 22'd2183985;
                12'd1995: exp <= 22'd2182378;
                12'd1996: exp <= 22'd2180771;
                12'd1997: exp <= 22'd2179163;
                12'd1998: exp <= 22'd2177556;
                12'd1999: exp <= 22'd2175949;
                12'd2000: exp <= 22'd2174341;
                12'd2001: exp <= 22'd2172734;
                12'd2002: exp <= 22'd2171126;
                12'd2003: exp <= 22'd2169519;
                12'd2004: exp <= 22'd2167911;
                12'd2005: exp <= 22'd2166304;
                12'd2006: exp <= 22'd2164696;
                12'd2007: exp <= 22'd2163088;
                12'd2008: exp <= 22'd2161481;
                12'd2009: exp <= 22'd2159873;
                12'd2010: exp <= 22'd2158265;
                12'd2011: exp <= 22'd2156657;
                12'd2012: exp <= 22'd2155049;
                12'd2013: exp <= 22'd2153442;
                12'd2014: exp <= 22'd2151834;
                12'd2015: exp <= 22'd2150226;
                12'd2016: exp <= 22'd2148618;
                12'd2017: exp <= 22'd2147010;
                12'd2018: exp <= 22'd2145402;
                12'd2019: exp <= 22'd2143794;
                12'd2020: exp <= 22'd2142185;
                12'd2021: exp <= 22'd2140577;
                12'd2022: exp <= 22'd2138969;
                12'd2023: exp <= 22'd2137361;
                12'd2024: exp <= 22'd2135753;
                12'd2025: exp <= 22'd2134144;
                12'd2026: exp <= 22'd2132536;
                12'd2027: exp <= 22'd2130928;
                12'd2028: exp <= 22'd2129320;
                12'd2029: exp <= 22'd2127711;
                12'd2030: exp <= 22'd2126103;
                12'd2031: exp <= 22'd2124495;
                12'd2032: exp <= 22'd2122886;
                12'd2033: exp <= 22'd2121278;
                12'd2034: exp <= 22'd2119670;
                12'd2035: exp <= 22'd2118061;
                12'd2036: exp <= 22'd2116453;
                12'd2037: exp <= 22'd2114844;
                12'd2038: exp <= 22'd2113236;
                12'd2039: exp <= 22'd2111627;
                12'd2040: exp <= 22'd2110019;
                12'd2041: exp <= 22'd2108410;
                12'd2042: exp <= 22'd2106802;
                12'd2043: exp <= 22'd2105193;
                12'd2044: exp <= 22'd2103585;
                12'd2045: exp <= 22'd2101976;
                12'd2046: exp <= 22'd2100368;
                12'd2047: exp <= 22'd2098759;
                12'd2048: exp <= 22'd2097151;
                12'd2049: exp <= 22'd2095543;
                12'd2050: exp <= 22'd2093934;
                12'd2051: exp <= 22'd2092326;
                12'd2052: exp <= 22'd2090717;
                12'd2053: exp <= 22'd2089109;
                12'd2054: exp <= 22'd2087500;
                12'd2055: exp <= 22'd2085892;
                12'd2056: exp <= 22'd2084283;
                12'd2057: exp <= 22'd2082675;
                12'd2058: exp <= 22'd2081066;
                12'd2059: exp <= 22'd2079458;
                12'd2060: exp <= 22'd2077849;
                12'd2061: exp <= 22'd2076241;
                12'd2062: exp <= 22'd2074632;
                12'd2063: exp <= 22'd2073024;
                12'd2064: exp <= 22'd2071416;
                12'd2065: exp <= 22'd2069807;
                12'd2066: exp <= 22'd2068199;
                12'd2067: exp <= 22'd2066591;
                12'd2068: exp <= 22'd2064982;
                12'd2069: exp <= 22'd2063374;
                12'd2070: exp <= 22'd2061766;
                12'd2071: exp <= 22'd2060158;
                12'd2072: exp <= 22'd2058549;
                12'd2073: exp <= 22'd2056941;
                12'd2074: exp <= 22'd2055333;
                12'd2075: exp <= 22'd2053725;
                12'd2076: exp <= 22'd2052117;
                12'd2077: exp <= 22'd2050508;
                12'd2078: exp <= 22'd2048900;
                12'd2079: exp <= 22'd2047292;
                12'd2080: exp <= 22'd2045684;
                12'd2081: exp <= 22'd2044076;
                12'd2082: exp <= 22'd2042468;
                12'd2083: exp <= 22'd2040860;
                12'd2084: exp <= 22'd2039253;
                12'd2085: exp <= 22'd2037645;
                12'd2086: exp <= 22'd2036037;
                12'd2087: exp <= 22'd2034429;
                12'd2088: exp <= 22'd2032821;
                12'd2089: exp <= 22'd2031214;
                12'd2090: exp <= 22'd2029606;
                12'd2091: exp <= 22'd2027998;
                12'd2092: exp <= 22'd2026391;
                12'd2093: exp <= 22'd2024783;
                12'd2094: exp <= 22'd2023176;
                12'd2095: exp <= 22'd2021568;
                12'd2096: exp <= 22'd2019961;
                12'd2097: exp <= 22'd2018353;
                12'd2098: exp <= 22'd2016746;
                12'd2099: exp <= 22'd2015139;
                12'd2100: exp <= 22'd2013531;
                12'd2101: exp <= 22'd2011924;
                12'd2102: exp <= 22'd2010317;
                12'd2103: exp <= 22'd2008710;
                12'd2104: exp <= 22'd2007103;
                12'd2105: exp <= 22'd2005496;
                12'd2106: exp <= 22'd2003889;
                12'd2107: exp <= 22'd2002282;
                12'd2108: exp <= 22'd2000675;
                12'd2109: exp <= 22'd1999069;
                12'd2110: exp <= 22'd1997462;
                12'd2111: exp <= 22'd1995855;
                12'd2112: exp <= 22'd1994249;
                12'd2113: exp <= 22'd1992642;
                12'd2114: exp <= 22'd1991036;
                12'd2115: exp <= 22'd1989429;
                12'd2116: exp <= 22'd1987823;
                12'd2117: exp <= 22'd1986217;
                12'd2118: exp <= 22'd1984610;
                12'd2119: exp <= 22'd1983004;
                12'd2120: exp <= 22'd1981398;
                12'd2121: exp <= 22'd1979792;
                12'd2122: exp <= 22'd1978186;
                12'd2123: exp <= 22'd1976580;
                12'd2124: exp <= 22'd1974975;
                12'd2125: exp <= 22'd1973369;
                12'd2126: exp <= 22'd1971763;
                12'd2127: exp <= 22'd1970158;
                12'd2128: exp <= 22'd1968552;
                12'd2129: exp <= 22'd1966947;
                12'd2130: exp <= 22'd1965341;
                12'd2131: exp <= 22'd1963736;
                12'd2132: exp <= 22'd1962131;
                12'd2133: exp <= 22'd1960526;
                12'd2134: exp <= 22'd1958921;
                12'd2135: exp <= 22'd1957316;
                12'd2136: exp <= 22'd1955711;
                12'd2137: exp <= 22'd1954106;
                12'd2138: exp <= 22'd1952501;
                12'd2139: exp <= 22'd1950897;
                12'd2140: exp <= 22'd1949292;
                12'd2141: exp <= 22'd1947688;
                12'd2142: exp <= 22'd1946083;
                12'd2143: exp <= 22'd1944479;
                12'd2144: exp <= 22'd1942875;
                12'd2145: exp <= 22'd1941271;
                12'd2146: exp <= 22'd1939667;
                12'd2147: exp <= 22'd1938063;
                12'd2148: exp <= 22'd1936459;
                12'd2149: exp <= 22'd1934855;
                12'd2150: exp <= 22'd1933252;
                12'd2151: exp <= 22'd1931648;
                12'd2152: exp <= 22'd1930045;
                12'd2153: exp <= 22'd1928441;
                12'd2154: exp <= 22'd1926838;
                12'd2155: exp <= 22'd1925235;
                12'd2156: exp <= 22'd1923632;
                12'd2157: exp <= 22'd1922029;
                12'd2158: exp <= 22'd1920426;
                12'd2159: exp <= 22'd1918824;
                12'd2160: exp <= 22'd1917221;
                12'd2161: exp <= 22'd1915618;
                12'd2162: exp <= 22'd1914016;
                12'd2163: exp <= 22'd1912414;
                12'd2164: exp <= 22'd1910812;
                12'd2165: exp <= 22'd1909210;
                12'd2166: exp <= 22'd1907608;
                12'd2167: exp <= 22'd1906006;
                12'd2168: exp <= 22'd1904404;
                12'd2169: exp <= 22'd1902802;
                12'd2170: exp <= 22'd1901201;
                12'd2171: exp <= 22'd1899599;
                12'd2172: exp <= 22'd1897998;
                12'd2173: exp <= 22'd1896397;
                12'd2174: exp <= 22'd1894796;
                12'd2175: exp <= 22'd1893195;
                12'd2176: exp <= 22'd1891594;
                12'd2177: exp <= 22'd1889993;
                12'd2178: exp <= 22'd1888393;
                12'd2179: exp <= 22'd1886792;
                12'd2180: exp <= 22'd1885192;
                12'd2181: exp <= 22'd1883592;
                12'd2182: exp <= 22'd1881992;
                12'd2183: exp <= 22'd1880392;
                12'd2184: exp <= 22'd1878792;
                12'd2185: exp <= 22'd1877192;
                12'd2186: exp <= 22'd1875593;
                12'd2187: exp <= 22'd1873993;
                12'd2188: exp <= 22'd1872394;
                12'd2189: exp <= 22'd1870795;
                12'd2190: exp <= 22'd1869196;
                12'd2191: exp <= 22'd1867597;
                12'd2192: exp <= 22'd1865998;
                12'd2193: exp <= 22'd1864400;
                12'd2194: exp <= 22'd1862801;
                12'd2195: exp <= 22'd1861203;
                12'd2196: exp <= 22'd1859605;
                12'd2197: exp <= 22'd1858007;
                12'd2198: exp <= 22'd1856409;
                12'd2199: exp <= 22'd1854811;
                12'd2200: exp <= 22'd1853213;
                12'd2201: exp <= 22'd1851616;
                12'd2202: exp <= 22'd1850018;
                12'd2203: exp <= 22'd1848421;
                12'd2204: exp <= 22'd1846824;
                12'd2205: exp <= 22'd1845227;
                12'd2206: exp <= 22'd1843630;
                12'd2207: exp <= 22'd1842034;
                12'd2208: exp <= 22'd1840437;
                12'd2209: exp <= 22'd1838841;
                12'd2210: exp <= 22'd1837245;
                12'd2211: exp <= 22'd1835649;
                12'd2212: exp <= 22'd1834053;
                12'd2213: exp <= 22'd1832457;
                12'd2214: exp <= 22'd1830862;
                12'd2215: exp <= 22'd1829266;
                12'd2216: exp <= 22'd1827671;
                12'd2217: exp <= 22'd1826076;
                12'd2218: exp <= 22'd1824481;
                12'd2219: exp <= 22'd1822886;
                12'd2220: exp <= 22'd1821292;
                12'd2221: exp <= 22'd1819697;
                12'd2222: exp <= 22'd1818103;
                12'd2223: exp <= 22'd1816509;
                12'd2224: exp <= 22'd1814915;
                12'd2225: exp <= 22'd1813321;
                12'd2226: exp <= 22'd1811727;
                12'd2227: exp <= 22'd1810134;
                12'd2228: exp <= 22'd1808541;
                12'd2229: exp <= 22'd1806948;
                12'd2230: exp <= 22'd1805355;
                12'd2231: exp <= 22'd1803762;
                12'd2232: exp <= 22'd1802169;
                12'd2233: exp <= 22'd1800577;
                12'd2234: exp <= 22'd1798985;
                12'd2235: exp <= 22'd1797393;
                12'd2236: exp <= 22'd1795801;
                12'd2237: exp <= 22'd1794209;
                12'd2238: exp <= 22'd1792617;
                12'd2239: exp <= 22'd1791026;
                12'd2240: exp <= 22'd1789435;
                12'd2241: exp <= 22'd1787844;
                12'd2242: exp <= 22'd1786253;
                12'd2243: exp <= 22'd1784662;
                12'd2244: exp <= 22'd1783072;
                12'd2245: exp <= 22'd1781482;
                12'd2246: exp <= 22'd1779892;
                12'd2247: exp <= 22'd1778302;
                12'd2248: exp <= 22'd1776712;
                12'd2249: exp <= 22'd1775123;
                12'd2250: exp <= 22'd1773533;
                12'd2251: exp <= 22'd1771944;
                12'd2252: exp <= 22'd1770355;
                12'd2253: exp <= 22'd1768766;
                12'd2254: exp <= 22'd1767178;
                12'd2255: exp <= 22'd1765589;
                12'd2256: exp <= 22'd1764001;
                12'd2257: exp <= 22'd1762413;
                12'd2258: exp <= 22'd1760826;
                12'd2259: exp <= 22'd1759238;
                12'd2260: exp <= 22'd1757651;
                12'd2261: exp <= 22'd1756063;
                12'd2262: exp <= 22'd1754476;
                12'd2263: exp <= 22'd1752890;
                12'd2264: exp <= 22'd1751303;
                12'd2265: exp <= 22'd1749717;
                12'd2266: exp <= 22'd1748131;
                12'd2267: exp <= 22'd1746545;
                12'd2268: exp <= 22'd1744959;
                12'd2269: exp <= 22'd1743373;
                12'd2270: exp <= 22'd1741788;
                12'd2271: exp <= 22'd1740203;
                12'd2272: exp <= 22'd1738618;
                12'd2273: exp <= 22'd1737033;
                12'd2274: exp <= 22'd1735449;
                12'd2275: exp <= 22'd1733864;
                12'd2276: exp <= 22'd1732280;
                12'd2277: exp <= 22'd1730697;
                12'd2278: exp <= 22'd1729113;
                12'd2279: exp <= 22'd1727529;
                12'd2280: exp <= 22'd1725946;
                12'd2281: exp <= 22'd1724363;
                12'd2282: exp <= 22'd1722780;
                12'd2283: exp <= 22'd1721198;
                12'd2284: exp <= 22'd1719616;
                12'd2285: exp <= 22'd1718034;
                12'd2286: exp <= 22'd1716452;
                12'd2287: exp <= 22'd1714870;
                12'd2288: exp <= 22'd1713289;
                12'd2289: exp <= 22'd1711707;
                12'd2290: exp <= 22'd1710126;
                12'd2291: exp <= 22'd1708546;
                12'd2292: exp <= 22'd1706965;
                12'd2293: exp <= 22'd1705385;
                12'd2294: exp <= 22'd1703805;
                12'd2295: exp <= 22'd1702225;
                12'd2296: exp <= 22'd1700645;
                12'd2297: exp <= 22'd1699066;
                12'd2298: exp <= 22'd1697487;
                12'd2299: exp <= 22'd1695908;
                12'd2300: exp <= 22'd1694329;
                12'd2301: exp <= 22'd1692751;
                12'd2302: exp <= 22'd1691173;
                12'd2303: exp <= 22'd1689595;
                12'd2304: exp <= 22'd1688017;
                12'd2305: exp <= 22'd1686439;
                12'd2306: exp <= 22'd1684862;
                12'd2307: exp <= 22'd1683285;
                12'd2308: exp <= 22'd1681709;
                12'd2309: exp <= 22'd1680132;
                12'd2310: exp <= 22'd1678556;
                12'd2311: exp <= 22'd1676980;
                12'd2312: exp <= 22'd1675404;
                12'd2313: exp <= 22'd1673829;
                12'd2314: exp <= 22'd1672253;
                12'd2315: exp <= 22'd1670678;
                12'd2316: exp <= 22'd1669103;
                12'd2317: exp <= 22'd1667529;
                12'd2318: exp <= 22'd1665955;
                12'd2319: exp <= 22'd1664381;
                12'd2320: exp <= 22'd1662807;
                12'd2321: exp <= 22'd1661233;
                12'd2322: exp <= 22'd1659660;
                12'd2323: exp <= 22'd1658087;
                12'd2324: exp <= 22'd1656515;
                12'd2325: exp <= 22'd1654942;
                12'd2326: exp <= 22'd1653370;
                12'd2327: exp <= 22'd1651798;
                12'd2328: exp <= 22'd1650226;
                12'd2329: exp <= 22'd1648655;
                12'd2330: exp <= 22'd1647084;
                12'd2331: exp <= 22'd1645513;
                12'd2332: exp <= 22'd1643942;
                12'd2333: exp <= 22'd1642372;
                12'd2334: exp <= 22'd1640802;
                12'd2335: exp <= 22'd1639232;
                12'd2336: exp <= 22'd1637662;
                12'd2337: exp <= 22'd1636093;
                12'd2338: exp <= 22'd1634524;
                12'd2339: exp <= 22'd1632955;
                12'd2340: exp <= 22'd1631387;
                12'd2341: exp <= 22'd1629819;
                12'd2342: exp <= 22'd1628251;
                12'd2343: exp <= 22'd1626683;
                12'd2344: exp <= 22'd1625116;
                12'd2345: exp <= 22'd1623549;
                12'd2346: exp <= 22'd1621982;
                12'd2347: exp <= 22'd1620415;
                12'd2348: exp <= 22'd1618849;
                12'd2349: exp <= 22'd1617283;
                12'd2350: exp <= 22'd1615718;
                12'd2351: exp <= 22'd1614152;
                12'd2352: exp <= 22'd1612587;
                12'd2353: exp <= 22'd1611022;
                12'd2354: exp <= 22'd1609458;
                12'd2355: exp <= 22'd1607893;
                12'd2356: exp <= 22'd1606329;
                12'd2357: exp <= 22'd1604766;
                12'd2358: exp <= 22'd1603202;
                12'd2359: exp <= 22'd1601639;
                12'd2360: exp <= 22'd1600076;
                12'd2361: exp <= 22'd1598514;
                12'd2362: exp <= 22'd1596952;
                12'd2363: exp <= 22'd1595390;
                12'd2364: exp <= 22'd1593828;
                12'd2365: exp <= 22'd1592267;
                12'd2366: exp <= 22'd1590706;
                12'd2367: exp <= 22'd1589145;
                12'd2368: exp <= 22'd1587585;
                12'd2369: exp <= 22'd1586024;
                12'd2370: exp <= 22'd1584465;
                12'd2371: exp <= 22'd1582905;
                12'd2372: exp <= 22'd1581346;
                12'd2373: exp <= 22'd1579787;
                12'd2374: exp <= 22'd1578228;
                12'd2375: exp <= 22'd1576670;
                12'd2376: exp <= 22'd1575112;
                12'd2377: exp <= 22'd1573554;
                12'd2378: exp <= 22'd1571997;
                12'd2379: exp <= 22'd1570440;
                12'd2380: exp <= 22'd1568883;
                12'd2381: exp <= 22'd1567327;
                12'd2382: exp <= 22'd1565770;
                12'd2383: exp <= 22'd1564215;
                12'd2384: exp <= 22'd1562659;
                12'd2385: exp <= 22'd1561104;
                12'd2386: exp <= 22'd1559549;
                12'd2387: exp <= 22'd1557994;
                12'd2388: exp <= 22'd1556440;
                12'd2389: exp <= 22'd1554886;
                12'd2390: exp <= 22'd1553332;
                12'd2391: exp <= 22'd1551779;
                12'd2392: exp <= 22'd1550226;
                12'd2393: exp <= 22'd1548673;
                12'd2394: exp <= 22'd1547121;
                12'd2395: exp <= 22'd1545569;
                12'd2396: exp <= 22'd1544017;
                12'd2397: exp <= 22'd1542466;
                12'd2398: exp <= 22'd1540915;
                12'd2399: exp <= 22'd1539364;
                12'd2400: exp <= 22'd1537814;
                12'd2401: exp <= 22'd1536264;
                12'd2402: exp <= 22'd1534714;
                12'd2403: exp <= 22'd1533165;
                12'd2404: exp <= 22'd1531616;
                12'd2405: exp <= 22'd1530067;
                12'd2406: exp <= 22'd1528518;
                12'd2407: exp <= 22'd1526970;
                12'd2408: exp <= 22'd1525423;
                12'd2409: exp <= 22'd1523875;
                12'd2410: exp <= 22'd1522328;
                12'd2411: exp <= 22'd1520781;
                12'd2412: exp <= 22'd1519235;
                12'd2413: exp <= 22'd1517689;
                12'd2414: exp <= 22'd1516143;
                12'd2415: exp <= 22'd1514598;
                12'd2416: exp <= 22'd1513053;
                12'd2417: exp <= 22'd1511508;
                12'd2418: exp <= 22'd1509964;
                12'd2419: exp <= 22'd1508420;
                12'd2420: exp <= 22'd1506876;
                12'd2421: exp <= 22'd1505333;
                12'd2422: exp <= 22'd1503790;
                12'd2423: exp <= 22'd1502247;
                12'd2424: exp <= 22'd1500705;
                12'd2425: exp <= 22'd1499163;
                12'd2426: exp <= 22'd1497622;
                12'd2427: exp <= 22'd1496081;
                12'd2428: exp <= 22'd1494540;
                12'd2429: exp <= 22'd1492999;
                12'd2430: exp <= 22'd1491459;
                12'd2431: exp <= 22'd1489919;
                12'd2432: exp <= 22'd1488380;
                12'd2433: exp <= 22'd1486841;
                12'd2434: exp <= 22'd1485302;
                12'd2435: exp <= 22'd1483764;
                12'd2436: exp <= 22'd1482226;
                12'd2437: exp <= 22'd1480688;
                12'd2438: exp <= 22'd1479151;
                12'd2439: exp <= 22'd1477614;
                12'd2440: exp <= 22'd1476078;
                12'd2441: exp <= 22'd1474541;
                12'd2442: exp <= 22'd1473006;
                12'd2443: exp <= 22'd1471470;
                12'd2444: exp <= 22'd1469935;
                12'd2445: exp <= 22'd1468400;
                12'd2446: exp <= 22'd1466866;
                12'd2447: exp <= 22'd1465332;
                12'd2448: exp <= 22'd1463799;
                12'd2449: exp <= 22'd1462265;
                12'd2450: exp <= 22'd1460733;
                12'd2451: exp <= 22'd1459200;
                12'd2452: exp <= 22'd1457668;
                12'd2453: exp <= 22'd1456136;
                12'd2454: exp <= 22'd1454605;
                12'd2455: exp <= 22'd1453074;
                12'd2456: exp <= 22'd1451544;
                12'd2457: exp <= 22'd1450013;
                12'd2458: exp <= 22'd1448484;
                12'd2459: exp <= 22'd1446954;
                12'd2460: exp <= 22'd1445425;
                12'd2461: exp <= 22'd1443896;
                12'd2462: exp <= 22'd1442368;
                12'd2463: exp <= 22'd1440840;
                12'd2464: exp <= 22'd1439313;
                12'd2465: exp <= 22'd1437786;
                12'd2466: exp <= 22'd1436259;
                12'd2467: exp <= 22'd1434733;
                12'd2468: exp <= 22'd1433207;
                12'd2469: exp <= 22'd1431681;
                12'd2470: exp <= 22'd1430156;
                12'd2471: exp <= 22'd1428631;
                12'd2472: exp <= 22'd1427107;
                12'd2473: exp <= 22'd1425583;
                12'd2474: exp <= 22'd1424059;
                12'd2475: exp <= 22'd1422536;
                12'd2476: exp <= 22'd1421013;
                12'd2477: exp <= 22'd1419491;
                12'd2478: exp <= 22'd1417969;
                12'd2479: exp <= 22'd1416447;
                12'd2480: exp <= 22'd1414926;
                12'd2481: exp <= 22'd1413405;
                12'd2482: exp <= 22'd1411885;
                12'd2483: exp <= 22'd1410365;
                12'd2484: exp <= 22'd1408845;
                12'd2485: exp <= 22'd1407326;
                12'd2486: exp <= 22'd1405807;
                12'd2487: exp <= 22'd1404289;
                12'd2488: exp <= 22'd1402771;
                12'd2489: exp <= 22'd1401253;
                12'd2490: exp <= 22'd1399736;
                12'd2491: exp <= 22'd1398219;
                12'd2492: exp <= 22'd1396703;
                12'd2493: exp <= 22'd1395187;
                12'd2494: exp <= 22'd1393672;
                12'd2495: exp <= 22'd1392156;
                12'd2496: exp <= 22'd1390642;
                12'd2497: exp <= 22'd1389128;
                12'd2498: exp <= 22'd1387614;
                12'd2499: exp <= 22'd1386100;
                12'd2500: exp <= 22'd1384587;
                12'd2501: exp <= 22'd1383075;
                12'd2502: exp <= 22'd1381562;
                12'd2503: exp <= 22'd1380051;
                12'd2504: exp <= 22'd1378539;
                12'd2505: exp <= 22'd1377028;
                12'd2506: exp <= 22'd1375518;
                12'd2507: exp <= 22'd1374008;
                12'd2508: exp <= 22'd1372498;
                12'd2509: exp <= 22'd1370989;
                12'd2510: exp <= 22'd1369480;
                12'd2511: exp <= 22'd1367972;
                12'd2512: exp <= 22'd1366464;
                12'd2513: exp <= 22'd1364957;
                12'd2514: exp <= 22'd1363450;
                12'd2515: exp <= 22'd1361943;
                12'd2516: exp <= 22'd1360437;
                12'd2517: exp <= 22'd1358931;
                12'd2518: exp <= 22'd1357426;
                12'd2519: exp <= 22'd1355921;
                12'd2520: exp <= 22'd1354416;
                12'd2521: exp <= 22'd1352912;
                12'd2522: exp <= 22'd1351409;
                12'd2523: exp <= 22'd1349906;
                12'd2524: exp <= 22'd1348403;
                12'd2525: exp <= 22'd1346901;
                12'd2526: exp <= 22'd1345399;
                12'd2527: exp <= 22'd1343897;
                12'd2528: exp <= 22'd1342396;
                12'd2529: exp <= 22'd1340896;
                12'd2530: exp <= 22'd1339396;
                12'd2531: exp <= 22'd1337896;
                12'd2532: exp <= 22'd1336397;
                12'd2533: exp <= 22'd1334898;
                12'd2534: exp <= 22'd1333400;
                12'd2535: exp <= 22'd1331902;
                12'd2536: exp <= 22'd1330405;
                12'd2537: exp <= 22'd1328908;
                12'd2538: exp <= 22'd1327412;
                12'd2539: exp <= 22'd1325916;
                12'd2540: exp <= 22'd1324420;
                12'd2541: exp <= 22'd1322925;
                12'd2542: exp <= 22'd1321430;
                12'd2543: exp <= 22'd1319936;
                12'd2544: exp <= 22'd1318442;
                12'd2545: exp <= 22'd1316949;
                12'd2546: exp <= 22'd1315456;
                12'd2547: exp <= 22'd1313964;
                12'd2548: exp <= 22'd1312472;
                12'd2549: exp <= 22'd1310981;
                12'd2550: exp <= 22'd1309490;
                12'd2551: exp <= 22'd1307999;
                12'd2552: exp <= 22'd1306509;
                12'd2553: exp <= 22'd1305020;
                12'd2554: exp <= 22'd1303530;
                12'd2555: exp <= 22'd1302042;
                12'd2556: exp <= 22'd1300554;
                12'd2557: exp <= 22'd1299066;
                12'd2558: exp <= 22'd1297579;
                12'd2559: exp <= 22'd1296092;
                12'd2560: exp <= 22'd1294606;
                12'd2561: exp <= 22'd1293120;
                12'd2562: exp <= 22'd1291635;
                12'd2563: exp <= 22'd1290150;
                12'd2564: exp <= 22'd1288665;
                12'd2565: exp <= 22'd1287181;
                12'd2566: exp <= 22'd1285698;
                12'd2567: exp <= 22'd1284215;
                12'd2568: exp <= 22'd1282732;
                12'd2569: exp <= 22'd1281250;
                12'd2570: exp <= 22'd1279769;
                12'd2571: exp <= 22'd1278288;
                12'd2572: exp <= 22'd1276807;
                12'd2573: exp <= 22'd1275327;
                12'd2574: exp <= 22'd1273848;
                12'd2575: exp <= 22'd1272368;
                12'd2576: exp <= 22'd1270890;
                12'd2577: exp <= 22'd1269412;
                12'd2578: exp <= 22'd1267934;
                12'd2579: exp <= 22'd1266457;
                12'd2580: exp <= 22'd1264980;
                12'd2581: exp <= 22'd1263504;
                12'd2582: exp <= 22'd1262028;
                12'd2583: exp <= 22'd1260553;
                12'd2584: exp <= 22'd1259078;
                12'd2585: exp <= 22'd1257604;
                12'd2586: exp <= 22'd1256130;
                12'd2587: exp <= 22'd1254657;
                12'd2588: exp <= 22'd1253184;
                12'd2589: exp <= 22'd1251712;
                12'd2590: exp <= 22'd1250240;
                12'd2591: exp <= 22'd1248769;
                12'd2592: exp <= 22'd1247298;
                12'd2593: exp <= 22'd1245828;
                12'd2594: exp <= 22'd1244358;
                12'd2595: exp <= 22'd1242889;
                12'd2596: exp <= 22'd1241420;
                12'd2597: exp <= 22'd1239952;
                12'd2598: exp <= 22'd1238484;
                12'd2599: exp <= 22'd1237017;
                12'd2600: exp <= 22'd1235550;
                12'd2601: exp <= 22'd1234084;
                12'd2602: exp <= 22'd1232618;
                12'd2603: exp <= 22'd1231153;
                12'd2604: exp <= 22'd1229689;
                12'd2605: exp <= 22'd1228224;
                12'd2606: exp <= 22'd1226761;
                12'd2607: exp <= 22'd1225298;
                12'd2608: exp <= 22'd1223835;
                12'd2609: exp <= 22'd1222373;
                12'd2610: exp <= 22'd1220911;
                12'd2611: exp <= 22'd1219450;
                12'd2612: exp <= 22'd1217989;
                12'd2613: exp <= 22'd1216529;
                12'd2614: exp <= 22'd1215070;
                12'd2615: exp <= 22'd1213611;
                12'd2616: exp <= 22'd1212152;
                12'd2617: exp <= 22'd1210694;
                12'd2618: exp <= 22'd1209237;
                12'd2619: exp <= 22'd1207780;
                12'd2620: exp <= 22'd1206323;
                12'd2621: exp <= 22'd1204868;
                12'd2622: exp <= 22'd1203412;
                12'd2623: exp <= 22'd1201957;
                12'd2624: exp <= 22'd1200503;
                12'd2625: exp <= 22'd1199049;
                12'd2626: exp <= 22'd1197596;
                12'd2627: exp <= 22'd1196143;
                12'd2628: exp <= 22'd1194691;
                12'd2629: exp <= 22'd1193239;
                12'd2630: exp <= 22'd1191788;
                12'd2631: exp <= 22'd1190338;
                12'd2632: exp <= 22'd1188887;
                12'd2633: exp <= 22'd1187438;
                12'd2634: exp <= 22'd1185989;
                12'd2635: exp <= 22'd1184540;
                12'd2636: exp <= 22'd1183092;
                12'd2637: exp <= 22'd1181645;
                12'd2638: exp <= 22'd1180198;
                12'd2639: exp <= 22'd1178752;
                12'd2640: exp <= 22'd1177306;
                12'd2641: exp <= 22'd1175861;
                12'd2642: exp <= 22'd1174416;
                12'd2643: exp <= 22'd1172972;
                12'd2644: exp <= 22'd1171528;
                12'd2645: exp <= 22'd1170085;
                12'd2646: exp <= 22'd1168643;
                12'd2647: exp <= 22'd1167201;
                12'd2648: exp <= 22'd1165759;
                12'd2649: exp <= 22'd1164318;
                12'd2650: exp <= 22'd1162878;
                12'd2651: exp <= 22'd1161438;
                12'd2652: exp <= 22'd1159999;
                12'd2653: exp <= 22'd1158560;
                12'd2654: exp <= 22'd1157122;
                12'd2655: exp <= 22'd1155685;
                12'd2656: exp <= 22'd1154248;
                12'd2657: exp <= 22'd1152811;
                12'd2658: exp <= 22'd1151375;
                12'd2659: exp <= 22'd1149940;
                12'd2660: exp <= 22'd1148505;
                12'd2661: exp <= 22'd1147071;
                12'd2662: exp <= 22'd1145637;
                12'd2663: exp <= 22'd1144204;
                12'd2664: exp <= 22'd1142772;
                12'd2665: exp <= 22'd1141340;
                12'd2666: exp <= 22'd1139908;
                12'd2667: exp <= 22'd1138477;
                12'd2668: exp <= 22'd1137047;
                12'd2669: exp <= 22'd1135617;
                12'd2670: exp <= 22'd1134188;
                12'd2671: exp <= 22'd1132759;
                12'd2672: exp <= 22'd1131331;
                12'd2673: exp <= 22'd1129904;
                12'd2674: exp <= 22'd1128477;
                12'd2675: exp <= 22'd1127051;
                12'd2676: exp <= 22'd1125625;
                12'd2677: exp <= 22'd1124200;
                12'd2678: exp <= 22'd1122775;
                12'd2679: exp <= 22'd1121351;
                12'd2680: exp <= 22'd1119927;
                12'd2681: exp <= 22'd1118505;
                12'd2682: exp <= 22'd1117082;
                12'd2683: exp <= 22'd1115660;
                12'd2684: exp <= 22'd1114239;
                12'd2685: exp <= 22'd1112819;
                12'd2686: exp <= 22'd1111399;
                12'd2687: exp <= 22'd1109979;
                12'd2688: exp <= 22'd1108560;
                12'd2689: exp <= 22'd1107142;
                12'd2690: exp <= 22'd1105724;
                12'd2691: exp <= 22'd1104307;
                12'd2692: exp <= 22'd1102891;
                12'd2693: exp <= 22'd1101475;
                12'd2694: exp <= 22'd1100059;
                12'd2695: exp <= 22'd1098645;
                12'd2696: exp <= 22'd1097231;
                12'd2697: exp <= 22'd1095817;
                12'd2698: exp <= 22'd1094404;
                12'd2699: exp <= 22'd1092992;
                12'd2700: exp <= 22'd1091580;
                12'd2701: exp <= 22'd1090168;
                12'd2702: exp <= 22'd1088758;
                12'd2703: exp <= 22'd1087348;
                12'd2704: exp <= 22'd1085938;
                12'd2705: exp <= 22'd1084529;
                12'd2706: exp <= 22'd1083121;
                12'd2707: exp <= 22'd1081714;
                12'd2708: exp <= 22'd1080306;
                12'd2709: exp <= 22'd1078900;
                12'd2710: exp <= 22'd1077494;
                12'd2711: exp <= 22'd1076089;
                12'd2712: exp <= 22'd1074684;
                12'd2713: exp <= 22'd1073280;
                12'd2714: exp <= 22'd1071877;
                12'd2715: exp <= 22'd1070474;
                12'd2716: exp <= 22'd1069072;
                12'd2717: exp <= 22'd1067670;
                12'd2718: exp <= 22'd1066269;
                12'd2719: exp <= 22'd1064868;
                12'd2720: exp <= 22'd1063469;
                12'd2721: exp <= 22'd1062069;
                12'd2722: exp <= 22'd1060671;
                12'd2723: exp <= 22'd1059273;
                12'd2724: exp <= 22'd1057875;
                12'd2725: exp <= 22'd1056479;
                12'd2726: exp <= 22'd1055082;
                12'd2727: exp <= 22'd1053687;
                12'd2728: exp <= 22'd1052292;
                12'd2729: exp <= 22'd1050898;
                12'd2730: exp <= 22'd1049504;
                12'd2731: exp <= 22'd1048111;
                12'd2732: exp <= 22'd1046718;
                12'd2733: exp <= 22'd1045326;
                12'd2734: exp <= 22'd1043935;
                12'd2735: exp <= 22'd1042544;
                12'd2736: exp <= 22'd1041154;
                12'd2737: exp <= 22'd1039765;
                12'd2738: exp <= 22'd1038376;
                12'd2739: exp <= 22'd1036988;
                12'd2740: exp <= 22'd1035601;
                12'd2741: exp <= 22'd1034214;
                12'd2742: exp <= 22'd1032828;
                12'd2743: exp <= 22'd1031442;
                12'd2744: exp <= 22'd1030057;
                12'd2745: exp <= 22'd1028672;
                12'd2746: exp <= 22'd1027289;
                12'd2747: exp <= 22'd1025906;
                12'd2748: exp <= 22'd1024523;
                12'd2749: exp <= 22'd1023141;
                12'd2750: exp <= 22'd1021760;
                12'd2751: exp <= 22'd1020379;
                12'd2752: exp <= 22'd1018999;
                12'd2753: exp <= 22'd1017620;
                12'd2754: exp <= 22'd1016241;
                12'd2755: exp <= 22'd1014863;
                12'd2756: exp <= 22'd1013486;
                12'd2757: exp <= 22'd1012109;
                12'd2758: exp <= 22'd1010733;
                12'd2759: exp <= 22'd1009357;
                12'd2760: exp <= 22'd1007983;
                12'd2761: exp <= 22'd1006608;
                12'd2762: exp <= 22'd1005235;
                12'd2763: exp <= 22'd1003862;
                12'd2764: exp <= 22'd1002489;
                12'd2765: exp <= 22'd1001118;
                12'd2766: exp <= 22'd0999747;
                12'd2767: exp <= 22'd0998376;
                12'd2768: exp <= 22'd0997007;
                12'd2769: exp <= 22'd0995638;
                12'd2770: exp <= 22'd0994269;
                12'd2771: exp <= 22'd0992901;
                12'd2772: exp <= 22'd0991534;
                12'd2773: exp <= 22'd0990168;
                12'd2774: exp <= 22'd0988802;
                12'd2775: exp <= 22'd0987437;
                12'd2776: exp <= 22'd0986072;
                12'd2777: exp <= 22'd0984708;
                12'd2778: exp <= 22'd0983345;
                12'd2779: exp <= 22'd0981983;
                12'd2780: exp <= 22'd0980621;
                12'd2781: exp <= 22'd0979259;
                12'd2782: exp <= 22'd0977899;
                12'd2783: exp <= 22'd0976539;
                12'd2784: exp <= 22'd0975180;
                12'd2785: exp <= 22'd0973821;
                12'd2786: exp <= 22'd0972463;
                12'd2787: exp <= 22'd0971106;
                12'd2788: exp <= 22'd0969749;
                12'd2789: exp <= 22'd0968393;
                12'd2790: exp <= 22'd0967038;
                12'd2791: exp <= 22'd0965683;
                12'd2792: exp <= 22'd0964329;
                12'd2793: exp <= 22'd0962976;
                12'd2794: exp <= 22'd0961623;
                12'd2795: exp <= 22'd0960271;
                12'd2796: exp <= 22'd0958920;
                12'd2797: exp <= 22'd0957569;
                12'd2798: exp <= 22'd0956220;
                12'd2799: exp <= 22'd0954870;
                12'd2800: exp <= 22'd0953522;
                12'd2801: exp <= 22'd0952174;
                12'd2802: exp <= 22'd0950826;
                12'd2803: exp <= 22'd0949480;
                12'd2804: exp <= 22'd0948134;
                12'd2805: exp <= 22'd0946789;
                12'd2806: exp <= 22'd0945444;
                12'd2807: exp <= 22'd0944100;
                12'd2808: exp <= 22'd0942757;
                12'd2809: exp <= 22'd0941414;
                12'd2810: exp <= 22'd0940073;
                12'd2811: exp <= 22'd0938731;
                12'd2812: exp <= 22'd0937391;
                12'd2813: exp <= 22'd0936051;
                12'd2814: exp <= 22'd0934712;
                12'd2815: exp <= 22'd0933374;
                12'd2816: exp <= 22'd0932036;
                12'd2817: exp <= 22'd0930699;
                12'd2818: exp <= 22'd0929362;
                12'd2819: exp <= 22'd0928027;
                12'd2820: exp <= 22'd0926692;
                12'd2821: exp <= 22'd0925357;
                12'd2822: exp <= 22'd0924024;
                12'd2823: exp <= 22'd0922691;
                12'd2824: exp <= 22'd0921358;
                12'd2825: exp <= 22'd0920027;
                12'd2826: exp <= 22'd0918696;
                12'd2827: exp <= 22'd0917366;
                12'd2828: exp <= 22'd0916036;
                12'd2829: exp <= 22'd0914708;
                12'd2830: exp <= 22'd0913379;
                12'd2831: exp <= 22'd0912052;
                12'd2832: exp <= 22'd0910725;
                12'd2833: exp <= 22'd0909399;
                12'd2834: exp <= 22'd0908074;
                12'd2835: exp <= 22'd0906750;
                12'd2836: exp <= 22'd0905426;
                12'd2837: exp <= 22'd0904102;
                12'd2838: exp <= 22'd0902780;
                12'd2839: exp <= 22'd0901458;
                12'd2840: exp <= 22'd0900137;
                12'd2841: exp <= 22'd0898817;
                12'd2842: exp <= 22'd0897497;
                12'd2843: exp <= 22'd0896178;
                12'd2844: exp <= 22'd0894860;
                12'd2845: exp <= 22'd0893542;
                12'd2846: exp <= 22'd0892225;
                12'd2847: exp <= 22'd0890909;
                12'd2848: exp <= 22'd0889594;
                12'd2849: exp <= 22'd0888279;
                12'd2850: exp <= 22'd0886965;
                12'd2851: exp <= 22'd0885652;
                12'd2852: exp <= 22'd0884339;
                12'd2853: exp <= 22'd0883027;
                12'd2854: exp <= 22'd0881716;
                12'd2855: exp <= 22'd0880406;
                12'd2856: exp <= 22'd0879096;
                12'd2857: exp <= 22'd0877787;
                12'd2858: exp <= 22'd0876479;
                12'd2859: exp <= 22'd0875171;
                12'd2860: exp <= 22'd0873864;
                12'd2861: exp <= 22'd0872558;
                12'd2862: exp <= 22'd0871253;
                12'd2863: exp <= 22'd0869948;
                12'd2864: exp <= 22'd0868644;
                12'd2865: exp <= 22'd0867341;
                12'd2866: exp <= 22'd0866038;
                12'd2867: exp <= 22'd0864736;
                12'd2868: exp <= 22'd0863435;
                12'd2869: exp <= 22'd0862135;
                12'd2870: exp <= 22'd0860835;
                12'd2871: exp <= 22'd0859536;
                12'd2872: exp <= 22'd0858238;
                12'd2873: exp <= 22'd0856941;
                12'd2874: exp <= 22'd0855644;
                12'd2875: exp <= 22'd0854348;
                12'd2876: exp <= 22'd0853053;
                12'd2877: exp <= 22'd0851758;
                12'd2878: exp <= 22'd0850464;
                12'd2879: exp <= 22'd0849171;
                12'd2880: exp <= 22'd0847879;
                12'd2881: exp <= 22'd0846587;
                12'd2882: exp <= 22'd0845297;
                12'd2883: exp <= 22'd0844006;
                12'd2884: exp <= 22'd0842717;
                12'd2885: exp <= 22'd0841428;
                12'd2886: exp <= 22'd0840141;
                12'd2887: exp <= 22'd0838853;
                12'd2888: exp <= 22'd0837567;
                12'd2889: exp <= 22'd0836281;
                12'd2890: exp <= 22'd0834996;
                12'd2891: exp <= 22'd0833712;
                12'd2892: exp <= 22'd0832429;
                12'd2893: exp <= 22'd0831146;
                12'd2894: exp <= 22'd0829864;
                12'd2895: exp <= 22'd0828583;
                12'd2896: exp <= 22'd0827302;
                12'd2897: exp <= 22'd0826023;
                12'd2898: exp <= 22'd0824744;
                12'd2899: exp <= 22'd0823465;
                12'd2900: exp <= 22'd0822188;
                12'd2901: exp <= 22'd0820911;
                12'd2902: exp <= 22'd0819635;
                12'd2903: exp <= 22'd0818360;
                12'd2904: exp <= 22'd0817085;
                12'd2905: exp <= 22'd0815812;
                12'd2906: exp <= 22'd0814539;
                12'd2907: exp <= 22'd0813267;
                12'd2908: exp <= 22'd0811995;
                12'd2909: exp <= 22'd0810724;
                12'd2910: exp <= 22'd0809454;
                12'd2911: exp <= 22'd0808185;
                12'd2912: exp <= 22'd0806917;
                12'd2913: exp <= 22'd0805649;
                12'd2914: exp <= 22'd0804382;
                12'd2915: exp <= 22'd0803116;
                12'd2916: exp <= 22'd0801851;
                12'd2917: exp <= 22'd0800586;
                12'd2918: exp <= 22'd0799322;
                12'd2919: exp <= 22'd0798059;
                12'd2920: exp <= 22'd0796797;
                12'd2921: exp <= 22'd0795535;
                12'd2922: exp <= 22'd0794274;
                12'd2923: exp <= 22'd0793014;
                12'd2924: exp <= 22'd0791755;
                12'd2925: exp <= 22'd0790497;
                12'd2926: exp <= 22'd0789239;
                12'd2927: exp <= 22'd0787982;
                12'd2928: exp <= 22'd0786726;
                12'd2929: exp <= 22'd0785470;
                12'd2930: exp <= 22'd0784216;
                12'd2931: exp <= 22'd0782962;
                12'd2932: exp <= 22'd0781709;
                12'd2933: exp <= 22'd0780456;
                12'd2934: exp <= 22'd0779205;
                12'd2935: exp <= 22'd0777954;
                12'd2936: exp <= 22'd0776704;
                12'd2937: exp <= 22'd0775455;
                12'd2938: exp <= 22'd0774206;
                12'd2939: exp <= 22'd0772959;
                12'd2940: exp <= 22'd0771712;
                12'd2941: exp <= 22'd0770466;
                12'd2942: exp <= 22'd0769220;
                12'd2943: exp <= 22'd0767976;
                12'd2944: exp <= 22'd0766732;
                12'd2945: exp <= 22'd0765489;
                12'd2946: exp <= 22'd0764247;
                12'd2947: exp <= 22'd0763005;
                12'd2948: exp <= 22'd0761765;
                12'd2949: exp <= 22'd0760525;
                12'd2950: exp <= 22'd0759286;
                12'd2951: exp <= 22'd0758047;
                12'd2952: exp <= 22'd0756810;
                12'd2953: exp <= 22'd0755573;
                12'd2954: exp <= 22'd0754337;
                12'd2955: exp <= 22'd0753102;
                12'd2956: exp <= 22'd0751868;
                12'd2957: exp <= 22'd0750634;
                12'd2958: exp <= 22'd0749402;
                12'd2959: exp <= 22'd0748170;
                12'd2960: exp <= 22'd0746938;
                12'd2961: exp <= 22'd0745708;
                12'd2962: exp <= 22'd0744478;
                12'd2963: exp <= 22'd0743250;
                12'd2964: exp <= 22'd0742022;
                12'd2965: exp <= 22'd0740794;
                12'd2966: exp <= 22'd0739568;
                12'd2967: exp <= 22'd0738343;
                12'd2968: exp <= 22'd0737118;
                12'd2969: exp <= 22'd0735894;
                12'd2970: exp <= 22'd0734671;
                12'd2971: exp <= 22'd0733448;
                12'd2972: exp <= 22'd0732227;
                12'd2973: exp <= 22'd0731006;
                12'd2974: exp <= 22'd0729786;
                12'd2975: exp <= 22'd0728567;
                12'd2976: exp <= 22'd0727348;
                12'd2977: exp <= 22'd0726131;
                12'd2978: exp <= 22'd0724914;
                12'd2979: exp <= 22'd0723698;
                12'd2980: exp <= 22'd0722483;
                12'd2981: exp <= 22'd0721269;
                12'd2982: exp <= 22'd0720055;
                12'd2983: exp <= 22'd0718842;
                12'd2984: exp <= 22'd0717630;
                12'd2985: exp <= 22'd0716419;
                12'd2986: exp <= 22'd0715209;
                12'd2987: exp <= 22'd0714000;
                12'd2988: exp <= 22'd0712791;
                12'd2989: exp <= 22'd0711583;
                12'd2990: exp <= 22'd0710376;
                12'd2991: exp <= 22'd0709170;
                12'd2992: exp <= 22'd0707964;
                12'd2993: exp <= 22'd0706760;
                12'd2994: exp <= 22'd0705556;
                12'd2995: exp <= 22'd0704353;
                12'd2996: exp <= 22'd0703151;
                12'd2997: exp <= 22'd0701950;
                12'd2998: exp <= 22'd0700749;
                12'd2999: exp <= 22'd0699550;
                12'd3000: exp <= 22'd0698351;
                12'd3001: exp <= 22'd0697153;
                12'd3002: exp <= 22'd0695956;
                12'd3003: exp <= 22'd0694759;
                12'd3004: exp <= 22'd0693564;
                12'd3005: exp <= 22'd0692369;
                12'd3006: exp <= 22'd0691175;
                12'd3007: exp <= 22'd0689982;
                12'd3008: exp <= 22'd0688790;
                12'd3009: exp <= 22'd0687598;
                12'd3010: exp <= 22'd0686408;
                12'd3011: exp <= 22'd0685218;
                12'd3012: exp <= 22'd0684029;
                12'd3013: exp <= 22'd0682841;
                12'd3014: exp <= 22'd0681654;
                12'd3015: exp <= 22'd0680467;
                12'd3016: exp <= 22'd0679282;
                12'd3017: exp <= 22'd0678097;
                12'd3018: exp <= 22'd0676913;
                12'd3019: exp <= 22'd0675730;
                12'd3020: exp <= 22'd0674548;
                12'd3021: exp <= 22'd0673366;
                12'd3022: exp <= 22'd0672186;
                12'd3023: exp <= 22'd0671006;
                12'd3024: exp <= 22'd0669827;
                12'd3025: exp <= 22'd0668649;
                12'd3026: exp <= 22'd0667472;
                12'd3027: exp <= 22'd0666296;
                12'd3028: exp <= 22'd0665120;
                12'd3029: exp <= 22'd0663945;
                12'd3030: exp <= 22'd0662772;
                12'd3031: exp <= 22'd0661599;
                12'd3032: exp <= 22'd0660426;
                12'd3033: exp <= 22'd0659255;
                12'd3034: exp <= 22'd0658085;
                12'd3035: exp <= 22'd0656915;
                12'd3036: exp <= 22'd0655746;
                12'd3037: exp <= 22'd0654578;
                12'd3038: exp <= 22'd0653411;
                12'd3039: exp <= 22'd0652245;
                12'd3040: exp <= 22'd0651080;
                12'd3041: exp <= 22'd0649915;
                12'd3042: exp <= 22'd0648751;
                12'd3043: exp <= 22'd0647589;
                12'd3044: exp <= 22'd0646427;
                12'd3045: exp <= 22'd0645266;
                12'd3046: exp <= 22'd0644105;
                12'd3047: exp <= 22'd0642946;
                12'd3048: exp <= 22'd0641787;
                12'd3049: exp <= 22'd0640630;
                12'd3050: exp <= 22'd0639473;
                12'd3051: exp <= 22'd0638317;
                12'd3052: exp <= 22'd0637162;
                12'd3053: exp <= 22'd0636007;
                12'd3054: exp <= 22'd0634854;
                12'd3055: exp <= 22'd0633702;
                12'd3056: exp <= 22'd0632550;
                12'd3057: exp <= 22'd0631399;
                12'd3058: exp <= 22'd0630249;
                12'd3059: exp <= 22'd0629100;
                12'd3060: exp <= 22'd0627952;
                12'd3061: exp <= 22'd0626804;
                12'd3062: exp <= 22'd0625658;
                12'd3063: exp <= 22'd0624512;
                12'd3064: exp <= 22'd0623367;
                12'd3065: exp <= 22'd0622224;
                12'd3066: exp <= 22'd0621081;
                12'd3067: exp <= 22'd0619938;
                12'd3068: exp <= 22'd0618797;
                12'd3069: exp <= 22'd0617657;
                12'd3070: exp <= 22'd0616517;
                12'd3071: exp <= 22'd0615378;
                12'd3072: exp <= 22'd0614241;
                12'd3073: exp <= 22'd0613104;
                12'd3074: exp <= 22'd0611968;
                12'd3075: exp <= 22'd0610832;
                12'd3076: exp <= 22'd0609698;
                12'd3077: exp <= 22'd0608565;
                12'd3078: exp <= 22'd0607432;
                12'd3079: exp <= 22'd0606300;
                12'd3080: exp <= 22'd0605170;
                12'd3081: exp <= 22'd0604040;
                12'd3082: exp <= 22'd0602911;
                12'd3083: exp <= 22'd0601782;
                12'd3084: exp <= 22'd0600655;
                12'd3085: exp <= 22'd0599529;
                12'd3086: exp <= 22'd0598403;
                12'd3087: exp <= 22'd0597278;
                12'd3088: exp <= 22'd0596155;
                12'd3089: exp <= 22'd0595032;
                12'd3090: exp <= 22'd0593910;
                12'd3091: exp <= 22'd0592789;
                12'd3092: exp <= 22'd0591668;
                12'd3093: exp <= 22'd0590549;
                12'd3094: exp <= 22'd0589431;
                12'd3095: exp <= 22'd0588313;
                12'd3096: exp <= 22'd0587196;
                12'd3097: exp <= 22'd0586080;
                12'd3098: exp <= 22'd0584966;
                12'd3099: exp <= 22'd0583852;
                12'd3100: exp <= 22'd0582738;
                12'd3101: exp <= 22'd0581626;
                12'd3102: exp <= 22'd0580515;
                12'd3103: exp <= 22'd0579404;
                12'd3104: exp <= 22'd0578295;
                12'd3105: exp <= 22'd0577186;
                12'd3106: exp <= 22'd0576078;
                12'd3107: exp <= 22'd0574971;
                12'd3108: exp <= 22'd0573865;
                12'd3109: exp <= 22'd0572760;
                12'd3110: exp <= 22'd0571656;
                12'd3111: exp <= 22'd0570553;
                12'd3112: exp <= 22'd0569450;
                12'd3113: exp <= 22'd0568349;
                12'd3114: exp <= 22'd0567248;
                12'd3115: exp <= 22'd0566149;
                12'd3116: exp <= 22'd0565050;
                12'd3117: exp <= 22'd0563952;
                12'd3118: exp <= 22'd0562855;
                12'd3119: exp <= 22'd0561759;
                12'd3120: exp <= 22'd0560664;
                12'd3121: exp <= 22'd0559569;
                12'd3122: exp <= 22'd0558476;
                12'd3123: exp <= 22'd0557383;
                12'd3124: exp <= 22'd0556292;
                12'd3125: exp <= 22'd0555201;
                12'd3126: exp <= 22'd0554111;
                12'd3127: exp <= 22'd0553023;
                12'd3128: exp <= 22'd0551935;
                12'd3129: exp <= 22'd0550848;
                12'd3130: exp <= 22'd0549761;
                12'd3131: exp <= 22'd0548676;
                12'd3132: exp <= 22'd0547592;
                12'd3133: exp <= 22'd0546509;
                12'd3134: exp <= 22'd0545426;
                12'd3135: exp <= 22'd0544345;
                12'd3136: exp <= 22'd0543264;
                12'd3137: exp <= 22'd0542184;
                12'd3138: exp <= 22'd0541105;
                12'd3139: exp <= 22'd0540027;
                12'd3140: exp <= 22'd0538950;
                12'd3141: exp <= 22'd0537874;
                12'd3142: exp <= 22'd0536799;
                12'd3143: exp <= 22'd0535725;
                12'd3144: exp <= 22'd0534652;
                12'd3145: exp <= 22'd0533579;
                12'd3146: exp <= 22'd0532508;
                12'd3147: exp <= 22'd0531437;
                12'd3148: exp <= 22'd0530367;
                12'd3149: exp <= 22'd0529299;
                12'd3150: exp <= 22'd0528231;
                12'd3151: exp <= 22'd0527164;
                12'd3152: exp <= 22'd0526098;
                12'd3153: exp <= 22'd0525033;
                12'd3154: exp <= 22'd0523969;
                12'd3155: exp <= 22'd0522906;
                12'd3156: exp <= 22'd0521844;
                12'd3157: exp <= 22'd0520782;
                12'd3158: exp <= 22'd0519722;
                12'd3159: exp <= 22'd0518662;
                12'd3160: exp <= 22'd0517604;
                12'd3161: exp <= 22'd0516546;
                12'd3162: exp <= 22'd0515489;
                12'd3163: exp <= 22'd0514434;
                12'd3164: exp <= 22'd0513379;
                12'd3165: exp <= 22'd0512325;
                12'd3166: exp <= 22'd0511272;
                12'd3167: exp <= 22'd0510220;
                12'd3168: exp <= 22'd0509169;
                12'd3169: exp <= 22'd0508119;
                12'd3170: exp <= 22'd0507070;
                12'd3171: exp <= 22'd0506021;
                12'd3172: exp <= 22'd0504974;
                12'd3173: exp <= 22'd0503928;
                12'd3174: exp <= 22'd0502882;
                12'd3175: exp <= 22'd0501837;
                12'd3176: exp <= 22'd0500794;
                12'd3177: exp <= 22'd0499751;
                12'd3178: exp <= 22'd0498710;
                12'd3179: exp <= 22'd0497669;
                12'd3180: exp <= 22'd0496629;
                12'd3181: exp <= 22'd0495590;
                12'd3182: exp <= 22'd0494552;
                12'd3183: exp <= 22'd0493515;
                12'd3184: exp <= 22'd0492479;
                12'd3185: exp <= 22'd0491444;
                12'd3186: exp <= 22'd0490410;
                12'd3187: exp <= 22'd0489376;
                12'd3188: exp <= 22'd0488344;
                12'd3189: exp <= 22'd0487313;
                12'd3190: exp <= 22'd0486282;
                12'd3191: exp <= 22'd0485253;
                12'd3192: exp <= 22'd0484224;
                12'd3193: exp <= 22'd0483197;
                12'd3194: exp <= 22'd0482170;
                12'd3195: exp <= 22'd0481145;
                12'd3196: exp <= 22'd0480120;
                12'd3197: exp <= 22'd0479096;
                12'd3198: exp <= 22'd0478073;
                12'd3199: exp <= 22'd0477051;
                12'd3200: exp <= 22'd0476031;
                12'd3201: exp <= 22'd0475011;
                12'd3202: exp <= 22'd0473992;
                12'd3203: exp <= 22'd0472974;
                12'd3204: exp <= 22'd0471957;
                12'd3205: exp <= 22'd0470940;
                12'd3206: exp <= 22'd0469925;
                12'd3207: exp <= 22'd0468911;
                12'd3208: exp <= 22'd0467898;
                12'd3209: exp <= 22'd0466886;
                12'd3210: exp <= 22'd0465874;
                12'd3211: exp <= 22'd0464864;
                12'd3212: exp <= 22'd0463854;
                12'd3213: exp <= 22'd0462846;
                12'd3214: exp <= 22'd0461838;
                12'd3215: exp <= 22'd0460832;
                12'd3216: exp <= 22'd0459826;
                12'd3217: exp <= 22'd0458822;
                12'd3218: exp <= 22'd0457818;
                12'd3219: exp <= 22'd0456815;
                12'd3220: exp <= 22'd0455814;
                12'd3221: exp <= 22'd0454813;
                12'd3222: exp <= 22'd0453813;
                12'd3223: exp <= 22'd0452814;
                12'd3224: exp <= 22'd0451817;
                12'd3225: exp <= 22'd0450820;
                12'd3226: exp <= 22'd0449824;
                12'd3227: exp <= 22'd0448829;
                12'd3228: exp <= 22'd0447835;
                12'd3229: exp <= 22'd0446842;
                12'd3230: exp <= 22'd0445850;
                12'd3231: exp <= 22'd0444859;
                12'd3232: exp <= 22'd0443869;
                12'd3233: exp <= 22'd0442880;
                12'd3234: exp <= 22'd0441891;
                12'd3235: exp <= 22'd0440904;
                12'd3236: exp <= 22'd0439918;
                12'd3237: exp <= 22'd0438933;
                12'd3238: exp <= 22'd0437949;
                12'd3239: exp <= 22'd0436965;
                12'd3240: exp <= 22'd0435983;
                12'd3241: exp <= 22'd0435002;
                12'd3242: exp <= 22'd0434021;
                12'd3243: exp <= 22'd0433042;
                12'd3244: exp <= 22'd0432064;
                12'd3245: exp <= 22'd0431086;
                12'd3246: exp <= 22'd0430110;
                12'd3247: exp <= 22'd0429134;
                12'd3248: exp <= 22'd0428160;
                12'd3249: exp <= 22'd0427187;
                12'd3250: exp <= 22'd0426214;
                12'd3251: exp <= 22'd0425243;
                12'd3252: exp <= 22'd0424272;
                12'd3253: exp <= 22'd0423303;
                12'd3254: exp <= 22'd0422334;
                12'd3255: exp <= 22'd0421366;
                12'd3256: exp <= 22'd0420400;
                12'd3257: exp <= 22'd0419434;
                12'd3258: exp <= 22'd0418470;
                12'd3259: exp <= 22'd0417506;
                12'd3260: exp <= 22'd0416543;
                12'd3261: exp <= 22'd0415582;
                12'd3262: exp <= 22'd0414621;
                12'd3263: exp <= 22'd0413661;
                12'd3264: exp <= 22'd0412703;
                12'd3265: exp <= 22'd0411745;
                12'd3266: exp <= 22'd0410788;
                12'd3267: exp <= 22'd0409833;
                12'd3268: exp <= 22'd0408878;
                12'd3269: exp <= 22'd0407924;
                12'd3270: exp <= 22'd0406971;
                12'd3271: exp <= 22'd0406020;
                12'd3272: exp <= 22'd0405069;
                12'd3273: exp <= 22'd0404119;
                12'd3274: exp <= 22'd0403171;
                12'd3275: exp <= 22'd0402223;
                12'd3276: exp <= 22'd0401276;
                12'd3277: exp <= 22'd0400330;
                12'd3278: exp <= 22'd0399386;
                12'd3279: exp <= 22'd0398442;
                12'd3280: exp <= 22'd0397499;
                12'd3281: exp <= 22'd0396557;
                12'd3282: exp <= 22'd0395617;
                12'd3283: exp <= 22'd0394677;
                12'd3284: exp <= 22'd0393738;
                12'd3285: exp <= 22'd0392800;
                12'd3286: exp <= 22'd0391864;
                12'd3287: exp <= 22'd0390928;
                12'd3288: exp <= 22'd0389993;
                12'd3289: exp <= 22'd0389059;
                12'd3290: exp <= 22'd0388127;
                12'd3291: exp <= 22'd0387195;
                12'd3292: exp <= 22'd0386264;
                12'd3293: exp <= 22'd0385334;
                12'd3294: exp <= 22'd0384406;
                12'd3295: exp <= 22'd0383478;
                12'd3296: exp <= 22'd0382551;
                12'd3297: exp <= 22'd0381626;
                12'd3298: exp <= 22'd0380701;
                12'd3299: exp <= 22'd0379777;
                12'd3300: exp <= 22'd0378855;
                12'd3301: exp <= 22'd0377933;
                12'd3302: exp <= 22'd0377012;
                12'd3303: exp <= 22'd0376093;
                12'd3304: exp <= 22'd0375174;
                12'd3305: exp <= 22'd0374257;
                12'd3306: exp <= 22'd0373340;
                12'd3307: exp <= 22'd0372424;
                12'd3308: exp <= 22'd0371510;
                12'd3309: exp <= 22'd0370596;
                12'd3310: exp <= 22'd0369684;
                12'd3311: exp <= 22'd0368772;
                12'd3312: exp <= 22'd0367862;
                12'd3313: exp <= 22'd0366952;
                12'd3314: exp <= 22'd0366044;
                12'd3315: exp <= 22'd0365137;
                12'd3316: exp <= 22'd0364230;
                12'd3317: exp <= 22'd0363325;
                12'd3318: exp <= 22'd0362420;
                12'd3319: exp <= 22'd0361517;
                12'd3320: exp <= 22'd0360615;
                12'd3321: exp <= 22'd0359713;
                12'd3322: exp <= 22'd0358813;
                12'd3323: exp <= 22'd0357914;
                12'd3324: exp <= 22'd0357016;
                12'd3325: exp <= 22'd0356118;
                12'd3326: exp <= 22'd0355222;
                12'd3327: exp <= 22'd0354327;
                12'd3328: exp <= 22'd0353433;
                12'd3329: exp <= 22'd0352540;
                12'd3330: exp <= 22'd0351648;
                12'd3331: exp <= 22'd0350757;
                12'd3332: exp <= 22'd0349867;
                12'd3333: exp <= 22'd0348978;
                12'd3334: exp <= 22'd0348090;
                12'd3335: exp <= 22'd0347203;
                12'd3336: exp <= 22'd0346317;
                12'd3337: exp <= 22'd0345432;
                12'd3338: exp <= 22'd0344548;
                12'd3339: exp <= 22'd0343665;
                12'd3340: exp <= 22'd0342783;
                12'd3341: exp <= 22'd0341902;
                12'd3342: exp <= 22'd0341023;
                12'd3343: exp <= 22'd0340144;
                12'd3344: exp <= 22'd0339266;
                12'd3345: exp <= 22'd0338390;
                12'd3346: exp <= 22'd0337514;
                12'd3347: exp <= 22'd0336640;
                12'd3348: exp <= 22'd0335766;
                12'd3349: exp <= 22'd0334894;
                12'd3350: exp <= 22'd0334022;
                12'd3351: exp <= 22'd0333152;
                12'd3352: exp <= 22'd0332282;
                12'd3353: exp <= 22'd0331414;
                12'd3354: exp <= 22'd0330547;
                12'd3355: exp <= 22'd0329680;
                12'd3356: exp <= 22'd0328815;
                12'd3357: exp <= 22'd0327951;
                12'd3358: exp <= 22'd0327088;
                12'd3359: exp <= 22'd0326226;
                12'd3360: exp <= 22'd0325365;
                12'd3361: exp <= 22'd0324505;
                12'd3362: exp <= 22'd0323646;
                12'd3363: exp <= 22'd0322788;
                12'd3364: exp <= 22'd0321931;
                12'd3365: exp <= 22'd0321075;
                12'd3366: exp <= 22'd0320220;
                12'd3367: exp <= 22'd0319366;
                12'd3368: exp <= 22'd0318514;
                12'd3369: exp <= 22'd0317662;
                12'd3370: exp <= 22'd0316811;
                12'd3371: exp <= 22'd0315962;
                12'd3372: exp <= 22'd0315113;
                12'd3373: exp <= 22'd0314266;
                12'd3374: exp <= 22'd0313419;
                12'd3375: exp <= 22'd0312574;
                12'd3376: exp <= 22'd0311730;
                12'd3377: exp <= 22'd0310886;
                12'd3378: exp <= 22'd0310044;
                12'd3379: exp <= 22'd0309203;
                12'd3380: exp <= 22'd0308363;
                12'd3381: exp <= 22'd0307524;
                12'd3382: exp <= 22'd0306686;
                12'd3383: exp <= 22'd0305849;
                12'd3384: exp <= 22'd0305013;
                12'd3385: exp <= 22'd0304178;
                12'd3386: exp <= 22'd0303344;
                12'd3387: exp <= 22'd0302512;
                12'd3388: exp <= 22'd0301680;
                12'd3389: exp <= 22'd0300849;
                12'd3390: exp <= 22'd0300020;
                12'd3391: exp <= 22'd0299191;
                12'd3392: exp <= 22'd0298364;
                12'd3393: exp <= 22'd0297537;
                12'd3394: exp <= 22'd0296712;
                12'd3395: exp <= 22'd0295888;
                12'd3396: exp <= 22'd0295064;
                12'd3397: exp <= 22'd0294242;
                12'd3398: exp <= 22'd0293421;
                12'd3399: exp <= 22'd0292601;
                12'd3400: exp <= 22'd0291782;
                12'd3401: exp <= 22'd0290964;
                12'd3402: exp <= 22'd0290147;
                12'd3403: exp <= 22'd0289332;
                12'd3404: exp <= 22'd0288517;
                12'd3405: exp <= 22'd0287703;
                12'd3406: exp <= 22'd0286891;
                12'd3407: exp <= 22'd0286079;
                12'd3408: exp <= 22'd0285269;
                12'd3409: exp <= 22'd0284459;
                12'd3410: exp <= 22'd0283651;
                12'd3411: exp <= 22'd0282844;
                12'd3412: exp <= 22'd0282037;
                12'd3413: exp <= 22'd0281232;
                12'd3414: exp <= 22'd0280428;
                12'd3415: exp <= 22'd0279625;
                12'd3416: exp <= 22'd0278823;
                12'd3417: exp <= 22'd0278022;
                12'd3418: exp <= 22'd0277223;
                12'd3419: exp <= 22'd0276424;
                12'd3420: exp <= 22'd0275626;
                12'd3421: exp <= 22'd0274830;
                12'd3422: exp <= 22'd0274034;
                12'd3423: exp <= 22'd0273240;
                12'd3424: exp <= 22'd0272446;
                12'd3425: exp <= 22'd0271654;
                12'd3426: exp <= 22'd0270863;
                12'd3427: exp <= 22'd0270073;
                12'd3428: exp <= 22'd0269284;
                12'd3429: exp <= 22'd0268496;
                12'd3430: exp <= 22'd0267709;
                12'd3431: exp <= 22'd0266923;
                12'd3432: exp <= 22'd0266138;
                12'd3433: exp <= 22'd0265354;
                12'd3434: exp <= 22'd0264572;
                12'd3435: exp <= 22'd0263790;
                12'd3436: exp <= 22'd0263010;
                12'd3437: exp <= 22'd0262230;
                12'd3438: exp <= 22'd0261452;
                12'd3439: exp <= 22'd0260675;
                12'd3440: exp <= 22'd0259899;
                12'd3441: exp <= 22'd0259124;
                12'd3442: exp <= 22'd0258350;
                12'd3443: exp <= 22'd0257577;
                12'd3444: exp <= 22'd0256805;
                12'd3445: exp <= 22'd0256034;
                12'd3446: exp <= 22'd0255265;
                12'd3447: exp <= 22'd0254496;
                12'd3448: exp <= 22'd0253729;
                12'd3449: exp <= 22'd0252962;
                12'd3450: exp <= 22'd0252197;
                12'd3451: exp <= 22'd0251433;
                12'd3452: exp <= 22'd0250670;
                12'd3453: exp <= 22'd0249908;
                12'd3454: exp <= 22'd0249147;
                12'd3455: exp <= 22'd0248387;
                12'd3456: exp <= 22'd0247628;
                12'd3457: exp <= 22'd0246870;
                12'd3458: exp <= 22'd0246114;
                12'd3459: exp <= 22'd0245358;
                12'd3460: exp <= 22'd0244604;
                12'd3461: exp <= 22'd0243850;
                12'd3462: exp <= 22'd0243098;
                12'd3463: exp <= 22'd0242347;
                12'd3464: exp <= 22'd0241597;
                12'd3465: exp <= 22'd0240848;
                12'd3466: exp <= 22'd0240100;
                12'd3467: exp <= 22'd0239353;
                12'd3468: exp <= 22'd0238608;
                12'd3469: exp <= 22'd0237863;
                12'd3470: exp <= 22'd0237120;
                12'd3471: exp <= 22'd0236377;
                12'd3472: exp <= 22'd0235636;
                12'd3473: exp <= 22'd0234896;
                12'd3474: exp <= 22'd0234156;
                12'd3475: exp <= 22'd0233418;
                12'd3476: exp <= 22'd0232681;
                12'd3477: exp <= 22'd0231946;
                12'd3478: exp <= 22'd0231211;
                12'd3479: exp <= 22'd0230477;
                12'd3480: exp <= 22'd0229745;
                12'd3481: exp <= 22'd0229013;
                12'd3482: exp <= 22'd0228283;
                12'd3483: exp <= 22'd0227554;
                12'd3484: exp <= 22'd0226825;
                12'd3485: exp <= 22'd0226098;
                12'd3486: exp <= 22'd0225372;
                12'd3487: exp <= 22'd0224648;
                12'd3488: exp <= 22'd0223924;
                12'd3489: exp <= 22'd0223201;
                12'd3490: exp <= 22'd0222480;
                12'd3491: exp <= 22'd0221759;
                12'd3492: exp <= 22'd0221040;
                12'd3493: exp <= 22'd0220322;
                12'd3494: exp <= 22'd0219605;
                12'd3495: exp <= 22'd0218889;
                12'd3496: exp <= 22'd0218174;
                12'd3497: exp <= 22'd0217460;
                12'd3498: exp <= 22'd0216747;
                12'd3499: exp <= 22'd0216035;
                12'd3500: exp <= 22'd0215325;
                12'd3501: exp <= 22'd0214616;
                12'd3502: exp <= 22'd0213907;
                12'd3503: exp <= 22'd0213200;
                12'd3504: exp <= 22'd0212494;
                12'd3505: exp <= 22'd0211789;
                12'd3506: exp <= 22'd0211085;
                12'd3507: exp <= 22'd0210383;
                12'd3508: exp <= 22'd0209681;
                12'd3509: exp <= 22'd0208980;
                12'd3510: exp <= 22'd0208281;
                12'd3511: exp <= 22'd0207583;
                12'd3512: exp <= 22'd0206885;
                12'd3513: exp <= 22'd0206189;
                12'd3514: exp <= 22'd0205494;
                12'd3515: exp <= 22'd0204801;
                12'd3516: exp <= 22'd0204108;
                12'd3517: exp <= 22'd0203416;
                12'd3518: exp <= 22'd0202726;
                12'd3519: exp <= 22'd0202036;
                12'd3520: exp <= 22'd0201348;
                12'd3521: exp <= 22'd0200661;
                12'd3522: exp <= 22'd0199975;
                12'd3523: exp <= 22'd0199290;
                12'd3524: exp <= 22'd0198606;
                12'd3525: exp <= 22'd0197923;
                12'd3526: exp <= 22'd0197242;
                12'd3527: exp <= 22'd0196561;
                12'd3528: exp <= 22'd0195882;
                12'd3529: exp <= 22'd0195204;
                12'd3530: exp <= 22'd0194527;
                12'd3531: exp <= 22'd0193851;
                12'd3532: exp <= 22'd0193176;
                12'd3533: exp <= 22'd0192502;
                12'd3534: exp <= 22'd0191829;
                12'd3535: exp <= 22'd0191158;
                12'd3536: exp <= 22'd0190488;
                12'd3537: exp <= 22'd0189818;
                12'd3538: exp <= 22'd0189150;
                12'd3539: exp <= 22'd0188483;
                12'd3540: exp <= 22'd0187817;
                12'd3541: exp <= 22'd0187152;
                12'd3542: exp <= 22'd0186489;
                12'd3543: exp <= 22'd0185826;
                12'd3544: exp <= 22'd0185165;
                12'd3545: exp <= 22'd0184505;
                12'd3546: exp <= 22'd0183845;
                12'd3547: exp <= 22'd0183187;
                12'd3548: exp <= 22'd0182531;
                12'd3549: exp <= 22'd0181875;
                12'd3550: exp <= 22'd0181220;
                12'd3551: exp <= 22'd0180567;
                12'd3552: exp <= 22'd0179914;
                12'd3553: exp <= 22'd0179263;
                12'd3554: exp <= 22'd0178613;
                12'd3555: exp <= 22'd0177964;
                12'd3556: exp <= 22'd0177316;
                12'd3557: exp <= 22'd0176669;
                12'd3558: exp <= 22'd0176024;
                12'd3559: exp <= 22'd0175379;
                12'd3560: exp <= 22'd0174736;
                12'd3561: exp <= 22'd0174093;
                12'd3562: exp <= 22'd0173452;
                12'd3563: exp <= 22'd0172812;
                12'd3564: exp <= 22'd0172174;
                12'd3565: exp <= 22'd0171536;
                12'd3566: exp <= 22'd0170899;
                12'd3567: exp <= 22'd0170264;
                12'd3568: exp <= 22'd0169630;
                12'd3569: exp <= 22'd0168996;
                12'd3570: exp <= 22'd0168364;
                12'd3571: exp <= 22'd0167733;
                12'd3572: exp <= 22'd0167104;
                12'd3573: exp <= 22'd0166475;
                12'd3574: exp <= 22'd0165848;
                12'd3575: exp <= 22'd0165221;
                12'd3576: exp <= 22'd0164596;
                12'd3577: exp <= 22'd0163972;
                12'd3578: exp <= 22'd0163349;
                12'd3579: exp <= 22'd0162727;
                12'd3580: exp <= 22'd0162106;
                12'd3581: exp <= 22'd0161487;
                12'd3582: exp <= 22'd0160869;
                12'd3583: exp <= 22'd0160251;
                12'd3584: exp <= 22'd0159635;
                12'd3585: exp <= 22'd0159020;
                12'd3586: exp <= 22'd0158406;
                12'd3587: exp <= 22'd0157794;
                12'd3588: exp <= 22'd0157182;
                12'd3589: exp <= 22'd0156572;
                12'd3590: exp <= 22'd0155962;
                12'd3591: exp <= 22'd0155354;
                12'd3592: exp <= 22'd0154747;
                12'd3593: exp <= 22'd0154141;
                12'd3594: exp <= 22'd0153537;
                12'd3595: exp <= 22'd0152933;
                12'd3596: exp <= 22'd0152331;
                12'd3597: exp <= 22'd0151730;
                12'd3598: exp <= 22'd0151129;
                12'd3599: exp <= 22'd0150530;
                12'd3600: exp <= 22'd0149933;
                12'd3601: exp <= 22'd0149336;
                12'd3602: exp <= 22'd0148740;
                12'd3603: exp <= 22'd0148146;
                12'd3604: exp <= 22'd0147553;
                12'd3605: exp <= 22'd0146961;
                12'd3606: exp <= 22'd0146370;
                12'd3607: exp <= 22'd0145780;
                12'd3608: exp <= 22'd0145191;
                12'd3609: exp <= 22'd0144604;
                12'd3610: exp <= 22'd0144017;
                12'd3611: exp <= 22'd0143432;
                12'd3612: exp <= 22'd0142848;
                12'd3613: exp <= 22'd0142265;
                12'd3614: exp <= 22'd0141683;
                12'd3615: exp <= 22'd0141103;
                12'd3616: exp <= 22'd0140523;
                12'd3617: exp <= 22'd0139945;
                12'd3618: exp <= 22'd0139368;
                12'd3619: exp <= 22'd0138792;
                12'd3620: exp <= 22'd0138217;
                12'd3621: exp <= 22'd0137643;
                12'd3622: exp <= 22'd0137071;
                12'd3623: exp <= 22'd0136499;
                12'd3624: exp <= 22'd0135929;
                12'd3625: exp <= 22'd0135360;
                12'd3626: exp <= 22'd0134792;
                12'd3627: exp <= 22'd0134225;
                12'd3628: exp <= 22'd0133660;
                12'd3629: exp <= 22'd0133095;
                12'd3630: exp <= 22'd0132532;
                12'd3631: exp <= 22'd0131970;
                12'd3632: exp <= 22'd0131409;
                12'd3633: exp <= 22'd0130849;
                12'd3634: exp <= 22'd0130290;
                12'd3635: exp <= 22'd0129733;
                12'd3636: exp <= 22'd0129176;
                12'd3637: exp <= 22'd0128621;
                12'd3638: exp <= 22'd0128067;
                12'd3639: exp <= 22'd0127514;
                12'd3640: exp <= 22'd0126962;
                12'd3641: exp <= 22'd0126412;
                12'd3642: exp <= 22'd0125862;
                12'd3643: exp <= 22'd0125314;
                12'd3644: exp <= 22'd0124767;
                12'd3645: exp <= 22'd0124221;
                12'd3646: exp <= 22'd0123676;
                12'd3647: exp <= 22'd0123132;
                12'd3648: exp <= 22'd0122590;
                12'd3649: exp <= 22'd0122049;
                12'd3650: exp <= 22'd0121509;
                12'd3651: exp <= 22'd0120970;
                12'd3652: exp <= 22'd0120432;
                12'd3653: exp <= 22'd0119895;
                12'd3654: exp <= 22'd0119360;
                12'd3655: exp <= 22'd0118825;
                12'd3656: exp <= 22'd0118292;
                12'd3657: exp <= 22'd0117760;
                12'd3658: exp <= 22'd0117229;
                12'd3659: exp <= 22'd0116700;
                12'd3660: exp <= 22'd0116171;
                12'd3661: exp <= 22'd0115644;
                12'd3662: exp <= 22'd0115118;
                12'd3663: exp <= 22'd0114593;
                12'd3664: exp <= 22'd0114069;
                12'd3665: exp <= 22'd0113546;
                12'd3666: exp <= 22'd0113025;
                12'd3667: exp <= 22'd0112504;
                12'd3668: exp <= 22'd0111985;
                12'd3669: exp <= 22'd0111467;
                12'd3670: exp <= 22'd0110950;
                12'd3671: exp <= 22'd0110434;
                12'd3672: exp <= 22'd0109920;
                12'd3673: exp <= 22'd0109407;
                12'd3674: exp <= 22'd0108894;
                12'd3675: exp <= 22'd0108383;
                12'd3676: exp <= 22'd0107874;
                12'd3677: exp <= 22'd0107365;
                12'd3678: exp <= 22'd0106858;
                12'd3679: exp <= 22'd0106351;
                12'd3680: exp <= 22'd0105846;
                12'd3681: exp <= 22'd0105342;
                12'd3682: exp <= 22'd0104839;
                12'd3683: exp <= 22'd0104338;
                12'd3684: exp <= 22'd0103837;
                12'd3685: exp <= 22'd0103338;
                12'd3686: exp <= 22'd0102840;
                12'd3687: exp <= 22'd0102343;
                12'd3688: exp <= 22'd0101847;
                12'd3689: exp <= 22'd0101353;
                12'd3690: exp <= 22'd0100859;
                12'd3691: exp <= 22'd0100367;
                12'd3692: exp <= 22'd0099876;
                12'd3693: exp <= 22'd0099386;
                12'd3694: exp <= 22'd0098897;
                12'd3695: exp <= 22'd0098410;
                12'd3696: exp <= 22'd0097923;
                12'd3697: exp <= 22'd0097438;
                12'd3698: exp <= 22'd0096954;
                12'd3699: exp <= 22'd0096471;
                12'd3700: exp <= 22'd0095990;
                12'd3701: exp <= 22'd0095509;
                12'd3702: exp <= 22'd0095030;
                12'd3703: exp <= 22'd0094552;
                12'd3704: exp <= 22'd0094075;
                12'd3705: exp <= 22'd0093599;
                12'd3706: exp <= 22'd0093124;
                12'd3707: exp <= 22'd0092651;
                12'd3708: exp <= 22'd0092179;
                12'd3709: exp <= 22'd0091708;
                12'd3710: exp <= 22'd0091238;
                12'd3711: exp <= 22'd0090769;
                12'd3712: exp <= 22'd0090302;
                12'd3713: exp <= 22'd0089835;
                12'd3714: exp <= 22'd0089370;
                12'd3715: exp <= 22'd0088906;
                12'd3716: exp <= 22'd0088443;
                12'd3717: exp <= 22'd0087982;
                12'd3718: exp <= 22'd0087521;
                12'd3719: exp <= 22'd0087062;
                12'd3720: exp <= 22'd0086604;
                12'd3721: exp <= 22'd0086147;
                12'd3722: exp <= 22'd0085692;
                12'd3723: exp <= 22'd0085237;
                12'd3724: exp <= 22'd0084784;
                12'd3725: exp <= 22'd0084332;
                12'd3726: exp <= 22'd0083881;
                12'd3727: exp <= 22'd0083431;
                12'd3728: exp <= 22'd0082982;
                12'd3729: exp <= 22'd0082535;
                12'd3730: exp <= 22'd0082089;
                12'd3731: exp <= 22'd0081644;
                12'd3732: exp <= 22'd0081200;
                12'd3733: exp <= 22'd0080757;
                12'd3734: exp <= 22'd0080316;
                12'd3735: exp <= 22'd0079875;
                12'd3736: exp <= 22'd0079436;
                12'd3737: exp <= 22'd0078998;
                12'd3738: exp <= 22'd0078562;
                12'd3739: exp <= 22'd0078126;
                12'd3740: exp <= 22'd0077692;
                12'd3741: exp <= 22'd0077258;
                12'd3742: exp <= 22'd0076826;
                12'd3743: exp <= 22'd0076396;
                12'd3744: exp <= 22'd0075966;
                12'd3745: exp <= 22'd0075538;
                12'd3746: exp <= 22'd0075110;
                12'd3747: exp <= 22'd0074684;
                12'd3748: exp <= 22'd0074260;
                12'd3749: exp <= 22'd0073836;
                12'd3750: exp <= 22'd0073413;
                12'd3751: exp <= 22'd0072992;
                12'd3752: exp <= 22'd0072572;
                12'd3753: exp <= 22'd0072153;
                12'd3754: exp <= 22'd0071736;
                12'd3755: exp <= 22'd0071319;
                12'd3756: exp <= 22'd0070904;
                12'd3757: exp <= 22'd0070490;
                12'd3758: exp <= 22'd0070077;
                12'd3759: exp <= 22'd0069665;
                12'd3760: exp <= 22'd0069254;
                12'd3761: exp <= 22'd0068845;
                12'd3762: exp <= 22'd0068437;
                12'd3763: exp <= 22'd0068030;
                12'd3764: exp <= 22'd0067624;
                12'd3765: exp <= 22'd0067220;
                12'd3766: exp <= 22'd0066816;
                12'd3767: exp <= 22'd0066414;
                12'd3768: exp <= 22'd0066013;
                12'd3769: exp <= 22'd0065613;
                12'd3770: exp <= 22'd0065215;
                12'd3771: exp <= 22'd0064817;
                12'd3772: exp <= 22'd0064421;
                12'd3773: exp <= 22'd0064026;
                12'd3774: exp <= 22'd0063632;
                12'd3775: exp <= 22'd0063239;
                12'd3776: exp <= 22'd0062848;
                12'd3777: exp <= 22'd0062458;
                12'd3778: exp <= 22'd0062069;
                12'd3779: exp <= 22'd0061681;
                12'd3780: exp <= 22'd0061294;
                12'd3781: exp <= 22'd0060909;
                12'd3782: exp <= 22'd0060525;
                12'd3783: exp <= 22'd0060142;
                12'd3784: exp <= 22'd0059760;
                12'd3785: exp <= 22'd0059379;
                12'd3786: exp <= 22'd0059000;
                12'd3787: exp <= 22'd0058621;
                12'd3788: exp <= 22'd0058244;
                12'd3789: exp <= 22'd0057868;
                12'd3790: exp <= 22'd0057494;
                12'd3791: exp <= 22'd0057120;
                12'd3792: exp <= 22'd0056748;
                12'd3793: exp <= 22'd0056377;
                12'd3794: exp <= 22'd0056007;
                12'd3795: exp <= 22'd0055638;
                12'd3796: exp <= 22'd0055271;
                12'd3797: exp <= 22'd0054905;
                12'd3798: exp <= 22'd0054540;
                12'd3799: exp <= 22'd0054176;
                12'd3800: exp <= 22'd0053813;
                12'd3801: exp <= 22'd0053452;
                12'd3802: exp <= 22'd0053092;
                12'd3803: exp <= 22'd0052732;
                12'd3804: exp <= 22'd0052375;
                12'd3805: exp <= 22'd0052018;
                12'd3806: exp <= 22'd0051663;
                12'd3807: exp <= 22'd0051308;
                12'd3808: exp <= 22'd0050955;
                12'd3809: exp <= 22'd0050604;
                12'd3810: exp <= 22'd0050253;
                12'd3811: exp <= 22'd0049903;
                12'd3812: exp <= 22'd0049555;
                12'd3813: exp <= 22'd0049208;
                12'd3814: exp <= 22'd0048862;
                12'd3815: exp <= 22'd0048518;
                12'd3816: exp <= 22'd0048174;
                12'd3817: exp <= 22'd0047832;
                12'd3818: exp <= 22'd0047491;
                12'd3819: exp <= 22'd0047152;
                12'd3820: exp <= 22'd0046813;
                12'd3821: exp <= 22'd0046476;
                12'd3822: exp <= 22'd0046139;
                12'd3823: exp <= 22'd0045805;
                12'd3824: exp <= 22'd0045471;
                12'd3825: exp <= 22'd0045138;
                12'd3826: exp <= 22'd0044807;
                12'd3827: exp <= 22'd0044477;
                12'd3828: exp <= 22'd0044148;
                12'd3829: exp <= 22'd0043820;
                12'd3830: exp <= 22'd0043494;
                12'd3831: exp <= 22'd0043168;
                12'd3832: exp <= 22'd0042844;
                12'd3833: exp <= 22'd0042521;
                12'd3834: exp <= 22'd0042200;
                12'd3835: exp <= 22'd0041879;
                12'd3836: exp <= 22'd0041560;
                12'd3837: exp <= 22'd0041242;
                12'd3838: exp <= 22'd0040925;
                12'd3839: exp <= 22'd0040610;
                12'd3840: exp <= 22'd0040295;
                12'd3841: exp <= 22'd0039982;
                12'd3842: exp <= 22'd0039670;
                12'd3843: exp <= 22'd0039359;
                12'd3844: exp <= 22'd0039050;
                12'd3845: exp <= 22'd0038741;
                12'd3846: exp <= 22'd0038434;
                12'd3847: exp <= 22'd0038128;
                12'd3848: exp <= 22'd0037824;
                12'd3849: exp <= 22'd0037520;
                12'd3850: exp <= 22'd0037218;
                12'd3851: exp <= 22'd0036917;
                12'd3852: exp <= 22'd0036617;
                12'd3853: exp <= 22'd0036318;
                12'd3854: exp <= 22'd0036021;
                12'd3855: exp <= 22'd0035724;
                12'd3856: exp <= 22'd0035429;
                12'd3857: exp <= 22'd0035136;
                12'd3858: exp <= 22'd0034843;
                12'd3859: exp <= 22'd0034552;
                12'd3860: exp <= 22'd0034261;
                12'd3861: exp <= 22'd0033972;
                12'd3862: exp <= 22'd0033685;
                12'd3863: exp <= 22'd0033398;
                12'd3864: exp <= 22'd0033113;
                12'd3865: exp <= 22'd0032829;
                12'd3866: exp <= 22'd0032546;
                12'd3867: exp <= 22'd0032264;
                12'd3868: exp <= 22'd0031984;
                12'd3869: exp <= 22'd0031704;
                12'd3870: exp <= 22'd0031426;
                12'd3871: exp <= 22'd0031150;
                12'd3872: exp <= 22'd0030874;
                12'd3873: exp <= 22'd0030600;
                12'd3874: exp <= 22'd0030326;
                12'd3875: exp <= 22'd0030055;
                12'd3876: exp <= 22'd0029784;
                12'd3877: exp <= 22'd0029514;
                12'd3878: exp <= 22'd0029246;
                12'd3879: exp <= 22'd0028979;
                12'd3880: exp <= 22'd0028713;
                12'd3881: exp <= 22'd0028448;
                12'd3882: exp <= 22'd0028185;
                12'd3883: exp <= 22'd0027923;
                12'd3884: exp <= 22'd0027662;
                12'd3885: exp <= 22'd0027402;
                12'd3886: exp <= 22'd0027143;
                12'd3887: exp <= 22'd0026886;
                12'd3888: exp <= 22'd0026630;
                12'd3889: exp <= 22'd0026375;
                12'd3890: exp <= 22'd0026121;
                12'd3891: exp <= 22'd0025869;
                12'd3892: exp <= 22'd0025618;
                12'd3893: exp <= 22'd0025367;
                12'd3894: exp <= 22'd0025119;
                12'd3895: exp <= 22'd0024871;
                12'd3896: exp <= 22'd0024625;
                12'd3897: exp <= 22'd0024380;
                12'd3898: exp <= 22'd0024136;
                12'd3899: exp <= 22'd0023893;
                12'd3900: exp <= 22'd0023651;
                12'd3901: exp <= 22'd0023411;
                12'd3902: exp <= 22'd0023172;
                12'd3903: exp <= 22'd0022934;
                12'd3904: exp <= 22'd0022698;
                12'd3905: exp <= 22'd0022462;
                12'd3906: exp <= 22'd0022228;
                12'd3907: exp <= 22'd0021995;
                12'd3908: exp <= 22'd0021763;
                12'd3909: exp <= 22'd0021533;
                12'd3910: exp <= 22'd0021303;
                12'd3911: exp <= 22'd0021075;
                12'd3912: exp <= 22'd0020848;
                12'd3913: exp <= 22'd0020623;
                12'd3914: exp <= 22'd0020398;
                12'd3915: exp <= 22'd0020175;
                12'd3916: exp <= 22'd0019953;
                12'd3917: exp <= 22'd0019732;
                12'd3918: exp <= 22'd0019513;
                12'd3919: exp <= 22'd0019295;
                12'd3920: exp <= 22'd0019078;
                12'd3921: exp <= 22'd0018862;
                12'd3922: exp <= 22'd0018647;
                12'd3923: exp <= 22'd0018434;
                12'd3924: exp <= 22'd0018221;
                12'd3925: exp <= 22'd0018010;
                12'd3926: exp <= 22'd0017801;
                12'd3927: exp <= 22'd0017592;
                12'd3928: exp <= 22'd0017385;
                12'd3929: exp <= 22'd0017179;
                12'd3930: exp <= 22'd0016974;
                12'd3931: exp <= 22'd0016770;
                12'd3932: exp <= 22'd0016568;
                12'd3933: exp <= 22'd0016367;
                12'd3934: exp <= 22'd0016167;
                12'd3935: exp <= 22'd0015968;
                12'd3936: exp <= 22'd0015771;
                12'd3937: exp <= 22'd0015574;
                12'd3938: exp <= 22'd0015379;
                12'd3939: exp <= 22'd0015185;
                12'd3940: exp <= 22'd0014993;
                12'd3941: exp <= 22'd0014801;
                12'd3942: exp <= 22'd0014611;
                12'd3943: exp <= 22'd0014422;
                12'd3944: exp <= 22'd0014235;
                12'd3945: exp <= 22'd0014048;
                12'd3946: exp <= 22'd0013863;
                12'd3947: exp <= 22'd0013679;
                12'd3948: exp <= 22'd0013496;
                12'd3949: exp <= 22'd0013314;
                12'd3950: exp <= 22'd0013134;
                12'd3951: exp <= 22'd0012955;
                12'd3952: exp <= 22'd0012777;
                12'd3953: exp <= 22'd0012600;
                12'd3954: exp <= 22'd0012425;
                12'd3955: exp <= 22'd0012251;
                12'd3956: exp <= 22'd0012078;
                12'd3957: exp <= 22'd0011906;
                12'd3958: exp <= 22'd0011735;
                12'd3959: exp <= 22'd0011566;
                12'd3960: exp <= 22'd0011398;
                12'd3961: exp <= 22'd0011231;
                12'd3962: exp <= 22'd0011065;
                12'd3963: exp <= 22'd0010901;
                12'd3964: exp <= 22'd0010738;
                12'd3965: exp <= 22'd0010576;
                12'd3966: exp <= 22'd0010415;
                12'd3967: exp <= 22'd0010256;
                12'd3968: exp <= 22'd0010097;
                12'd3969: exp <= 22'd0009940;
                12'd3970: exp <= 22'd0009784;
                12'd3971: exp <= 22'd0009630;
                12'd3972: exp <= 22'd0009477;
                12'd3973: exp <= 22'd0009324;
                12'd3974: exp <= 22'd0009174;
                12'd3975: exp <= 22'd0009024;
                12'd3976: exp <= 22'd0008875;
                12'd3977: exp <= 22'd0008728;
                12'd3978: exp <= 22'd0008582;
                12'd3979: exp <= 22'd0008437;
                12'd3980: exp <= 22'd0008294;
                12'd3981: exp <= 22'd0008152;
                12'd3982: exp <= 22'd0008010;
                12'd3983: exp <= 22'd0007871;
                12'd3984: exp <= 22'd0007732;
                12'd3985: exp <= 22'd0007595;
                12'd3986: exp <= 22'd0007458;
                12'd3987: exp <= 22'd0007324;
                12'd3988: exp <= 22'd0007190;
                12'd3989: exp <= 22'd0007057;
                12'd3990: exp <= 22'd0006926;
                12'd3991: exp <= 22'd0006796;
                12'd3992: exp <= 22'd0006667;
                12'd3993: exp <= 22'd0006540;
                12'd3994: exp <= 22'd0006413;
                12'd3995: exp <= 22'd0006288;
                12'd3996: exp <= 22'd0006164;
                12'd3997: exp <= 22'd0006042;
                12'd3998: exp <= 22'd0005920;
                12'd3999: exp <= 22'd0005800;
                12'd4000: exp <= 22'd0005681;
                12'd4001: exp <= 22'd0005564;
                12'd4002: exp <= 22'd0005447;
                12'd4003: exp <= 22'd0005332;
                12'd4004: exp <= 22'd0005218;
                12'd4005: exp <= 22'd0005105;
                12'd4006: exp <= 22'd0004994;
                12'd4007: exp <= 22'd0004883;
                12'd4008: exp <= 22'd0004774;
                12'd4009: exp <= 22'd0004666;
                12'd4010: exp <= 22'd0004560;
                12'd4011: exp <= 22'd0004454;
                12'd4012: exp <= 22'd0004350;
                12'd4013: exp <= 22'd0004247;
                12'd4014: exp <= 22'd0004145;
                12'd4015: exp <= 22'd0004045;
                12'd4016: exp <= 22'd0003946;
                12'd4017: exp <= 22'd0003848;
                12'd4018: exp <= 22'd0003751;
                12'd4019: exp <= 22'd0003655;
                12'd4020: exp <= 22'd0003561;
                12'd4021: exp <= 22'd0003468;
                12'd4022: exp <= 22'd0003376;
                12'd4023: exp <= 22'd0003285;
                12'd4024: exp <= 22'd0003196;
                12'd4025: exp <= 22'd0003108;
                12'd4026: exp <= 22'd0003021;
                12'd4027: exp <= 22'd0002935;
                12'd4028: exp <= 22'd0002851;
                12'd4029: exp <= 22'd0002767;
                12'd4030: exp <= 22'd0002685;
                12'd4031: exp <= 22'd0002605;
                12'd4032: exp <= 22'd0002525;
                12'd4033: exp <= 22'd0002447;
                12'd4034: exp <= 22'd0002370;
                12'd4035: exp <= 22'd0002294;
                12'd4036: exp <= 22'd0002219;
                12'd4037: exp <= 22'd0002146;
                12'd4038: exp <= 22'd0002074;
                12'd4039: exp <= 22'd0002003;
                12'd4040: exp <= 22'd0001933;
                12'd4041: exp <= 22'd0001865;
                12'd4042: exp <= 22'd0001797;
                12'd4043: exp <= 22'd0001731;
                12'd4044: exp <= 22'd0001667;
                12'd4045: exp <= 22'd0001603;
                12'd4046: exp <= 22'd0001541;
                12'd4047: exp <= 22'd0001480;
                12'd4048: exp <= 22'd0001420;
                12'd4049: exp <= 22'd0001361;
                12'd4050: exp <= 22'd0001304;
                12'd4051: exp <= 22'd0001248;
                12'd4052: exp <= 22'd0001193;
                12'd4053: exp <= 22'd0001139;
                12'd4054: exp <= 22'd0001087;
                12'd4055: exp <= 22'd0001036;
                12'd4056: exp <= 22'd0000986;
                12'd4057: exp <= 22'd0000937;
                12'd4058: exp <= 22'd0000890;
                12'd4059: exp <= 22'd0000843;
                12'd4060: exp <= 22'd0000798;
                12'd4061: exp <= 22'd0000755;
                12'd4062: exp <= 22'd0000712;
                12'd4063: exp <= 22'd0000671;
                12'd4064: exp <= 22'd0000631;
                12'd4065: exp <= 22'd0000592;
                12'd4066: exp <= 22'd0000554;
                12'd4067: exp <= 22'd0000518;
                12'd4068: exp <= 22'd0000483;
                12'd4069: exp <= 22'd0000449;
                12'd4070: exp <= 22'd0000416;
                12'd4071: exp <= 22'd0000385;
                12'd4072: exp <= 22'd0000354;
                12'd4073: exp <= 22'd0000325;
                12'd4074: exp <= 22'd0000298;
                12'd4075: exp <= 22'd0000271;
                12'd4076: exp <= 22'd0000246;
                12'd4077: exp <= 22'd0000222;
                12'd4078: exp <= 22'd0000199;
                12'd4079: exp <= 22'd0000177;
                12'd4080: exp <= 22'd0000157;
                12'd4081: exp <= 22'd0000138;
                12'd4082: exp <= 22'd0000120;
                12'd4083: exp <= 22'd0000103;
                12'd4084: exp <= 22'd0000088;
                12'd4085: exp <= 22'd0000074;
                12'd4086: exp <= 22'd0000061;
                12'd4087: exp <= 22'd0000049;
                12'd4088: exp <= 22'd0000038;
                12'd4089: exp <= 22'd0000029;
                12'd4090: exp <= 22'd0000021;
                12'd4091: exp <= 22'd0000014;
                12'd4092: exp <= 22'd0000009;
                12'd4093: exp <= 22'd0000005;
                12'd4094: exp <= 22'd0000001;
                12'd4095: exp <= 22'd0000000;
            endcase
        //2'b01: //linear
        //    exp = {addr, addr[19:18]};
    endcase
endmodule

/* This file is part of JT12 modification adding high precission audio
   mode called FM Overdrive

 
    JT12 program is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.

    JT12 program is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.

    You should have received a copy of the GNU General Public License
    along with JT12.  If not, see <http://www.gnu.org/licenses/>.

    Based on Sauraen VHDL version of OPN/OPN2, which is based on die shots.

    Author: Jose Tejada Gomez. Twitter: @topapate
    Version: 1.0
    Date: 27-1-2017 

*/

//altera message_off 10030

module jt12_logsin_hd
(
    input [15:0] addr,
    input clk, 
    input clk_en,
    input [1:0] fmo_sinelut,
    output reg [23:0] logsin
);

always @ (posedge clk) if(clk_en)
    case (fmo_sinelut)
        4'b00: //sinexp 12/24-bit
            case (addr[15:4])
                12'd0000: logsin <= 24'd00000000;
                12'd0001: logsin <= 24'd00000000;
                12'd0002: logsin <= 24'd00000001;
                12'd0003: logsin <= 24'd00000001;
                12'd0004: logsin <= 24'd00000002;
                12'd0005: logsin <= 24'd00000003;
                12'd0006: logsin <= 24'd00000005;
                12'd0007: logsin <= 24'd00000006;
                12'd0008: logsin <= 24'd00000008;
                12'd0009: logsin <= 24'd00000010;
                12'd0010: logsin <= 24'd00000012;
                12'd0011: logsin <= 24'd00000015;
                12'd0012: logsin <= 24'd00000017;
                12'd0013: logsin <= 24'd00000020;
                12'd0014: logsin <= 24'd00000023;
                12'd0015: logsin <= 24'd00000027;
                12'd0016: logsin <= 24'd00000030;
                12'd0017: logsin <= 24'd00000034;
                12'd0018: logsin <= 24'd00000038;
                12'd0019: logsin <= 24'd00000042;
                12'd0020: logsin <= 24'd00000047;
                12'd0021: logsin <= 24'd00000051;
                12'd0022: logsin <= 24'd00000056;
                12'd0023: logsin <= 24'd00000061;
                12'd0024: logsin <= 24'd00000067;
                12'd0025: logsin <= 24'd00000072;
                12'd0026: logsin <= 24'd00000078;
                12'd0027: logsin <= 24'd00000084;
                12'd0028: logsin <= 24'd00000090;
                12'd0029: logsin <= 24'd00000097;
                12'd0030: logsin <= 24'd00000103;
                12'd0031: logsin <= 24'd00000110;
                12'd0032: logsin <= 24'd00000118;
                12'd0033: logsin <= 24'd00000125;
                12'd0034: logsin <= 24'd00000132;
                12'd0035: logsin <= 24'd00000140;
                12'd0036: logsin <= 24'd00000148;
                12'd0037: logsin <= 24'd00000156;
                12'd0038: logsin <= 24'd00000165;
                12'd0039: logsin <= 24'd00000174;
                12'd0040: logsin <= 24'd00000182;
                12'd0041: logsin <= 24'd00000192;
                12'd0042: logsin <= 24'd00000201;
                12'd0043: logsin <= 24'd00000211;
                12'd0044: logsin <= 24'd00000220;
                12'd0045: logsin <= 24'd00000230;
                12'd0046: logsin <= 24'd00000241;
                12'd0047: logsin <= 24'd00000251;
                12'd0048: logsin <= 24'd00000262;
                12'd0049: logsin <= 24'd00000273;
                12'd0050: logsin <= 24'd00000284;
                12'd0051: logsin <= 24'd00000295;
                12'd0052: logsin <= 24'd00000307;
                12'd0053: logsin <= 24'd00000318;
                12'd0054: logsin <= 24'd00000330;
                12'd0055: logsin <= 24'd00000343;
                12'd0056: logsin <= 24'd00000355;
                12'd0057: logsin <= 24'd00000368;
                12'd0058: logsin <= 24'd00000381;
                12'd0059: logsin <= 24'd00000394;
                12'd0060: logsin <= 24'd00000407;
                12'd0061: logsin <= 24'd00000421;
                12'd0062: logsin <= 24'd00000435;
                12'd0063: logsin <= 24'd00000449;
                12'd0064: logsin <= 24'd00000463;
                12'd0065: logsin <= 24'd00000477;
                12'd0066: logsin <= 24'd00000492;
                12'd0067: logsin <= 24'd00000507;
                12'd0068: logsin <= 24'd00000522;
                12'd0069: logsin <= 24'd00000537;
                12'd0070: logsin <= 24'd00000553;
                12'd0071: logsin <= 24'd00000569;
                12'd0072: logsin <= 24'd00000585;
                12'd0073: logsin <= 24'd00000601;
                12'd0074: logsin <= 24'd00000617;
                12'd0075: logsin <= 24'd00000634;
                12'd0076: logsin <= 24'd00000651;
                12'd0077: logsin <= 24'd00000668;
                12'd0078: logsin <= 24'd00000686;
                12'd0079: logsin <= 24'd00000703;
                12'd0080: logsin <= 24'd00000721;
                12'd0081: logsin <= 24'd00000739;
                12'd0082: logsin <= 24'd00000757;
                12'd0083: logsin <= 24'd00000776;
                12'd0084: logsin <= 24'd00000794;
                12'd0085: logsin <= 24'd00000813;
                12'd0086: logsin <= 24'd00000832;
                12'd0087: logsin <= 24'd00000852;
                12'd0088: logsin <= 24'd00000871;
                12'd0089: logsin <= 24'd00000891;
                12'd0090: logsin <= 24'd00000911;
                12'd0091: logsin <= 24'd00000932;
                12'd0092: logsin <= 24'd00000952;
                12'd0093: logsin <= 24'd00000973;
                12'd0094: logsin <= 24'd00000994;
                12'd0095: logsin <= 24'd00001015;
                12'd0096: logsin <= 24'd00001036;
                12'd0097: logsin <= 24'd00001058;
                12'd0098: logsin <= 24'd00001080;
                12'd0099: logsin <= 24'd00001102;
                12'd0100: logsin <= 24'd00001124;
                12'd0101: logsin <= 24'd00001146;
                12'd0102: logsin <= 24'd00001169;
                12'd0103: logsin <= 24'd00001192;
                12'd0104: logsin <= 24'd00001215;
                12'd0105: logsin <= 24'd00001238;
                12'd0106: logsin <= 24'd00001262;
                12'd0107: logsin <= 24'd00001286;
                12'd0108: logsin <= 24'd00001310;
                12'd0109: logsin <= 24'd00001334;
                12'd0110: logsin <= 24'd00001359;
                12'd0111: logsin <= 24'd00001383;
                12'd0112: logsin <= 24'd00001408;
                12'd0113: logsin <= 24'd00001433;
                12'd0114: logsin <= 24'd00001459;
                12'd0115: logsin <= 24'd00001484;
                12'd0116: logsin <= 24'd00001510;
                12'd0117: logsin <= 24'd00001536;
                12'd0118: logsin <= 24'd00001563;
                12'd0119: logsin <= 24'd00001589;
                12'd0120: logsin <= 24'd00001616;
                12'd0121: logsin <= 24'd00001643;
                12'd0122: logsin <= 24'd00001670;
                12'd0123: logsin <= 24'd00001697;
                12'd0124: logsin <= 24'd00001725;
                12'd0125: logsin <= 24'd00001753;
                12'd0126: logsin <= 24'd00001781;
                12'd0127: logsin <= 24'd00001809;
                12'd0128: logsin <= 24'd00001838;
                12'd0129: logsin <= 24'd00001866;
                12'd0130: logsin <= 24'd00001895;
                12'd0131: logsin <= 24'd00001924;
                12'd0132: logsin <= 24'd00001954;
                12'd0133: logsin <= 24'd00001983;
                12'd0134: logsin <= 24'd00002013;
                12'd0135: logsin <= 24'd00002043;
                12'd0136: logsin <= 24'd00002074;
                12'd0137: logsin <= 24'd00002104;
                12'd0138: logsin <= 24'd00002135;
                12'd0139: logsin <= 24'd00002166;
                12'd0140: logsin <= 24'd00002197;
                12'd0141: logsin <= 24'd00002228;
                12'd0142: logsin <= 24'd00002260;
                12'd0143: logsin <= 24'd00002292;
                12'd0144: logsin <= 24'd00002324;
                12'd0145: logsin <= 24'd00002356;
                12'd0146: logsin <= 24'd00002389;
                12'd0147: logsin <= 24'd00002421;
                12'd0148: logsin <= 24'd00002454;
                12'd0149: logsin <= 24'd00002488;
                12'd0150: logsin <= 24'd00002521;
                12'd0151: logsin <= 24'd00002555;
                12'd0152: logsin <= 24'd00002589;
                12'd0153: logsin <= 24'd00002623;
                12'd0154: logsin <= 24'd00002657;
                12'd0155: logsin <= 24'd00002691;
                12'd0156: logsin <= 24'd00002726;
                12'd0157: logsin <= 24'd00002761;
                12'd0158: logsin <= 24'd00002796;
                12'd0159: logsin <= 24'd00002832;
                12'd0160: logsin <= 24'd00002867;
                12'd0161: logsin <= 24'd00002903;
                12'd0162: logsin <= 24'd00002939;
                12'd0163: logsin <= 24'd00002976;
                12'd0164: logsin <= 24'd00003012;
                12'd0165: logsin <= 24'd00003049;
                12'd0166: logsin <= 24'd00003086;
                12'd0167: logsin <= 24'd00003123;
                12'd0168: logsin <= 24'd00003161;
                12'd0169: logsin <= 24'd00003198;
                12'd0170: logsin <= 24'd00003236;
                12'd0171: logsin <= 24'd00003274;
                12'd0172: logsin <= 24'd00003313;
                12'd0173: logsin <= 24'd00003351;
                12'd0174: logsin <= 24'd00003390;
                12'd0175: logsin <= 24'd00003429;
                12'd0176: logsin <= 24'd00003468;
                12'd0177: logsin <= 24'd00003507;
                12'd0178: logsin <= 24'd00003547;
                12'd0179: logsin <= 24'd00003587;
                12'd0180: logsin <= 24'd00003627;
                12'd0181: logsin <= 24'd00003667;
                12'd0182: logsin <= 24'd00003708;
                12'd0183: logsin <= 24'd00003749;
                12'd0184: logsin <= 24'd00003790;
                12'd0185: logsin <= 24'd00003831;
                12'd0186: logsin <= 24'd00003873;
                12'd0187: logsin <= 24'd00003914;
                12'd0188: logsin <= 24'd00003956;
                12'd0189: logsin <= 24'd00003998;
                12'd0190: logsin <= 24'd00004041;
                12'd0191: logsin <= 24'd00004083;
                12'd0192: logsin <= 24'd00004126;
                12'd0193: logsin <= 24'd00004169;
                12'd0194: logsin <= 24'd00004212;
                12'd0195: logsin <= 24'd00004256;
                12'd0196: logsin <= 24'd00004299;
                12'd0197: logsin <= 24'd00004343;
                12'd0198: logsin <= 24'd00004387;
                12'd0199: logsin <= 24'd00004432;
                12'd0200: logsin <= 24'd00004476;
                12'd0201: logsin <= 24'd00004521;
                12'd0202: logsin <= 24'd00004566;
                12'd0203: logsin <= 24'd00004611;
                12'd0204: logsin <= 24'd00004657;
                12'd0205: logsin <= 24'd00004703;
                12'd0206: logsin <= 24'd00004749;
                12'd0207: logsin <= 24'd00004795;
                12'd0208: logsin <= 24'd00004841;
                12'd0209: logsin <= 24'd00004888;
                12'd0210: logsin <= 24'd00004934;
                12'd0211: logsin <= 24'd00004982;
                12'd0212: logsin <= 24'd00005029;
                12'd0213: logsin <= 24'd00005076;
                12'd0214: logsin <= 24'd00005124;
                12'd0215: logsin <= 24'd00005172;
                12'd0216: logsin <= 24'd00005220;
                12'd0217: logsin <= 24'd00005269;
                12'd0218: logsin <= 24'd00005317;
                12'd0219: logsin <= 24'd00005366;
                12'd0220: logsin <= 24'd00005415;
                12'd0221: logsin <= 24'd00005464;
                12'd0222: logsin <= 24'd00005514;
                12'd0223: logsin <= 24'd00005564;
                12'd0224: logsin <= 24'd00005614;
                12'd0225: logsin <= 24'd00005664;
                12'd0226: logsin <= 24'd00005714;
                12'd0227: logsin <= 24'd00005765;
                12'd0228: logsin <= 24'd00005816;
                12'd0229: logsin <= 24'd00005867;
                12'd0230: logsin <= 24'd00005918;
                12'd0231: logsin <= 24'd00005969;
                12'd0232: logsin <= 24'd00006021;
                12'd0233: logsin <= 24'd00006073;
                12'd0234: logsin <= 24'd00006125;
                12'd0235: logsin <= 24'd00006178;
                12'd0236: logsin <= 24'd00006231;
                12'd0237: logsin <= 24'd00006283;
                12'd0238: logsin <= 24'd00006336;
                12'd0239: logsin <= 24'd00006390;
                12'd0240: logsin <= 24'd00006443;
                12'd0241: logsin <= 24'd00006497;
                12'd0242: logsin <= 24'd00006551;
                12'd0243: logsin <= 24'd00006605;
                12'd0244: logsin <= 24'd00006660;
                12'd0245: logsin <= 24'd00006714;
                12'd0246: logsin <= 24'd00006769;
                12'd0247: logsin <= 24'd00006824;
                12'd0248: logsin <= 24'd00006880;
                12'd0249: logsin <= 24'd00006935;
                12'd0250: logsin <= 24'd00006991;
                12'd0251: logsin <= 24'd00007047;
                12'd0252: logsin <= 24'd00007103;
                12'd0253: logsin <= 24'd00007160;
                12'd0254: logsin <= 24'd00007217;
                12'd0255: logsin <= 24'd00007273;
                12'd0256: logsin <= 24'd00007331;
                12'd0257: logsin <= 24'd00007388;
                12'd0258: logsin <= 24'd00007446;
                12'd0259: logsin <= 24'd00007503;
                12'd0260: logsin <= 24'd00007561;
                12'd0261: logsin <= 24'd00007620;
                12'd0262: logsin <= 24'd00007678;
                12'd0263: logsin <= 24'd00007737;
                12'd0264: logsin <= 24'd00007796;
                12'd0265: logsin <= 24'd00007855;
                12'd0266: logsin <= 24'd00007914;
                12'd0267: logsin <= 24'd00007974;
                12'd0268: logsin <= 24'd00008034;
                12'd0269: logsin <= 24'd00008094;
                12'd0270: logsin <= 24'd00008154;
                12'd0271: logsin <= 24'd00008215;
                12'd0272: logsin <= 24'd00008275;
                12'd0273: logsin <= 24'd00008336;
                12'd0274: logsin <= 24'd00008398;
                12'd0275: logsin <= 24'd00008459;
                12'd0276: logsin <= 24'd00008521;
                12'd0277: logsin <= 24'd00008582;
                12'd0278: logsin <= 24'd00008645;
                12'd0279: logsin <= 24'd00008707;
                12'd0280: logsin <= 24'd00008769;
                12'd0281: logsin <= 24'd00008832;
                12'd0282: logsin <= 24'd00008895;
                12'd0283: logsin <= 24'd00008958;
                12'd0284: logsin <= 24'd00009022;
                12'd0285: logsin <= 24'd00009085;
                12'd0286: logsin <= 24'd00009149;
                12'd0287: logsin <= 24'd00009213;
                12'd0288: logsin <= 24'd00009278;
                12'd0289: logsin <= 24'd00009342;
                12'd0290: logsin <= 24'd00009407;
                12'd0291: logsin <= 24'd00009472;
                12'd0292: logsin <= 24'd00009537;
                12'd0293: logsin <= 24'd00009603;
                12'd0294: logsin <= 24'd00009669;
                12'd0295: logsin <= 24'd00009734;
                12'd0296: logsin <= 24'd00009801;
                12'd0297: logsin <= 24'd00009867;
                12'd0298: logsin <= 24'd00009934;
                12'd0299: logsin <= 24'd00010000;
                12'd0300: logsin <= 24'd00010067;
                12'd0301: logsin <= 24'd00010135;
                12'd0302: logsin <= 24'd00010202;
                12'd0303: logsin <= 24'd00010270;
                12'd0304: logsin <= 24'd00010338;
                12'd0305: logsin <= 24'd00010406;
                12'd0306: logsin <= 24'd00010474;
                12'd0307: logsin <= 24'd00010543;
                12'd0308: logsin <= 24'd00010612;
                12'd0309: logsin <= 24'd00010681;
                12'd0310: logsin <= 24'd00010750;
                12'd0311: logsin <= 24'd00010820;
                12'd0312: logsin <= 24'd00010889;
                12'd0313: logsin <= 24'd00010959;
                12'd0314: logsin <= 24'd00011030;
                12'd0315: logsin <= 24'd00011100;
                12'd0316: logsin <= 24'd00011171;
                12'd0317: logsin <= 24'd00011242;
                12'd0318: logsin <= 24'd00011313;
                12'd0319: logsin <= 24'd00011384;
                12'd0320: logsin <= 24'd00011456;
                12'd0321: logsin <= 24'd00011527;
                12'd0322: logsin <= 24'd00011599;
                12'd0323: logsin <= 24'd00011672;
                12'd0324: logsin <= 24'd00011744;
                12'd0325: logsin <= 24'd00011817;
                12'd0326: logsin <= 24'd00011890;
                12'd0327: logsin <= 24'd00011963;
                12'd0328: logsin <= 24'd00012036;
                12'd0329: logsin <= 24'd00012110;
                12'd0330: logsin <= 24'd00012184;
                12'd0331: logsin <= 24'd00012258;
                12'd0332: logsin <= 24'd00012332;
                12'd0333: logsin <= 24'd00012406;
                12'd0334: logsin <= 24'd00012481;
                12'd0335: logsin <= 24'd00012556;
                12'd0336: logsin <= 24'd00012631;
                12'd0337: logsin <= 24'd00012707;
                12'd0338: logsin <= 24'd00012782;
                12'd0339: logsin <= 24'd00012858;
                12'd0340: logsin <= 24'd00012934;
                12'd0341: logsin <= 24'd00013010;
                12'd0342: logsin <= 24'd00013087;
                12'd0343: logsin <= 24'd00013164;
                12'd0344: logsin <= 24'd00013241;
                12'd0345: logsin <= 24'd00013318;
                12'd0346: logsin <= 24'd00013395;
                12'd0347: logsin <= 24'd00013473;
                12'd0348: logsin <= 24'd00013551;
                12'd0349: logsin <= 24'd00013629;
                12'd0350: logsin <= 24'd00013707;
                12'd0351: logsin <= 24'd00013786;
                12'd0352: logsin <= 24'd00013865;
                12'd0353: logsin <= 24'd00013944;
                12'd0354: logsin <= 24'd00014023;
                12'd0355: logsin <= 24'd00014102;
                12'd0356: logsin <= 24'd00014182;
                12'd0357: logsin <= 24'd00014262;
                12'd0358: logsin <= 24'd00014342;
                12'd0359: logsin <= 24'd00014423;
                12'd0360: logsin <= 24'd00014503;
                12'd0361: logsin <= 24'd00014584;
                12'd0362: logsin <= 24'd00014665;
                12'd0363: logsin <= 24'd00014746;
                12'd0364: logsin <= 24'd00014828;
                12'd0365: logsin <= 24'd00014910;
                12'd0366: logsin <= 24'd00014992;
                12'd0367: logsin <= 24'd00015074;
                12'd0368: logsin <= 24'd00015156;
                12'd0369: logsin <= 24'd00015239;
                12'd0370: logsin <= 24'd00015322;
                12'd0371: logsin <= 24'd00015405;
                12'd0372: logsin <= 24'd00015488;
                12'd0373: logsin <= 24'd00015572;
                12'd0374: logsin <= 24'd00015655;
                12'd0375: logsin <= 24'd00015739;
                12'd0376: logsin <= 24'd00015824;
                12'd0377: logsin <= 24'd00015908;
                12'd0378: logsin <= 24'd00015993;
                12'd0379: logsin <= 24'd00016078;
                12'd0380: logsin <= 24'd00016163;
                12'd0381: logsin <= 24'd00016248;
                12'd0382: logsin <= 24'd00016334;
                12'd0383: logsin <= 24'd00016420;
                12'd0384: logsin <= 24'd00016506;
                12'd0385: logsin <= 24'd00016592;
                12'd0386: logsin <= 24'd00016679;
                12'd0387: logsin <= 24'd00016765;
                12'd0388: logsin <= 24'd00016852;
                12'd0389: logsin <= 24'd00016940;
                12'd0390: logsin <= 24'd00017027;
                12'd0391: logsin <= 24'd00017115;
                12'd0392: logsin <= 24'd00017202;
                12'd0393: logsin <= 24'd00017291;
                12'd0394: logsin <= 24'd00017379;
                12'd0395: logsin <= 24'd00017467;
                12'd0396: logsin <= 24'd00017556;
                12'd0397: logsin <= 24'd00017645;
                12'd0398: logsin <= 24'd00017734;
                12'd0399: logsin <= 24'd00017824;
                12'd0400: logsin <= 24'd00017914;
                12'd0401: logsin <= 24'd00018004;
                12'd0402: logsin <= 24'd00018094;
                12'd0403: logsin <= 24'd00018184;
                12'd0404: logsin <= 24'd00018275;
                12'd0405: logsin <= 24'd00018366;
                12'd0406: logsin <= 24'd00018457;
                12'd0407: logsin <= 24'd00018548;
                12'd0408: logsin <= 24'd00018639;
                12'd0409: logsin <= 24'd00018731;
                12'd0410: logsin <= 24'd00018823;
                12'd0411: logsin <= 24'd00018915;
                12'd0412: logsin <= 24'd00019008;
                12'd0413: logsin <= 24'd00019100;
                12'd0414: logsin <= 24'd00019193;
                12'd0415: logsin <= 24'd00019286;
                12'd0416: logsin <= 24'd00019380;
                12'd0417: logsin <= 24'd00019473;
                12'd0418: logsin <= 24'd00019567;
                12'd0419: logsin <= 24'd00019661;
                12'd0420: logsin <= 24'd00019755;
                12'd0421: logsin <= 24'd00019850;
                12'd0422: logsin <= 24'd00019945;
                12'd0423: logsin <= 24'd00020040;
                12'd0424: logsin <= 24'd00020135;
                12'd0425: logsin <= 24'd00020230;
                12'd0426: logsin <= 24'd00020326;
                12'd0427: logsin <= 24'd00020422;
                12'd0428: logsin <= 24'd00020518;
                12'd0429: logsin <= 24'd00020614;
                12'd0430: logsin <= 24'd00020711;
                12'd0431: logsin <= 24'd00020807;
                12'd0432: logsin <= 24'd00020904;
                12'd0433: logsin <= 24'd00021002;
                12'd0434: logsin <= 24'd00021099;
                12'd0435: logsin <= 24'd00021197;
                12'd0436: logsin <= 24'd00021295;
                12'd0437: logsin <= 24'd00021393;
                12'd0438: logsin <= 24'd00021491;
                12'd0439: logsin <= 24'd00021590;
                12'd0440: logsin <= 24'd00021689;
                12'd0441: logsin <= 24'd00021788;
                12'd0442: logsin <= 24'd00021887;
                12'd0443: logsin <= 24'd00021987;
                12'd0444: logsin <= 24'd00022086;
                12'd0445: logsin <= 24'd00022186;
                12'd0446: logsin <= 24'd00022286;
                12'd0447: logsin <= 24'd00022387;
                12'd0448: logsin <= 24'd00022488;
                12'd0449: logsin <= 24'd00022588;
                12'd0450: logsin <= 24'd00022690;
                12'd0451: logsin <= 24'd00022791;
                12'd0452: logsin <= 24'd00022893;
                12'd0453: logsin <= 24'd00022994;
                12'd0454: logsin <= 24'd00023096;
                12'd0455: logsin <= 24'd00023199;
                12'd0456: logsin <= 24'd00023301;
                12'd0457: logsin <= 24'd00023404;
                12'd0458: logsin <= 24'd00023507;
                12'd0459: logsin <= 24'd00023610;
                12'd0460: logsin <= 24'd00023713;
                12'd0461: logsin <= 24'd00023817;
                12'd0462: logsin <= 24'd00023921;
                12'd0463: logsin <= 24'd00024025;
                12'd0464: logsin <= 24'd00024129;
                12'd0465: logsin <= 24'd00024234;
                12'd0466: logsin <= 24'd00024339;
                12'd0467: logsin <= 24'd00024444;
                12'd0468: logsin <= 24'd00024549;
                12'd0469: logsin <= 24'd00024654;
                12'd0470: logsin <= 24'd00024760;
                12'd0471: logsin <= 24'd00024866;
                12'd0472: logsin <= 24'd00024972;
                12'd0473: logsin <= 24'd00025079;
                12'd0474: logsin <= 24'd00025185;
                12'd0475: logsin <= 24'd00025292;
                12'd0476: logsin <= 24'd00025399;
                12'd0477: logsin <= 24'd00025507;
                12'd0478: logsin <= 24'd00025614;
                12'd0479: logsin <= 24'd00025722;
                12'd0480: logsin <= 24'd00025830;
                12'd0481: logsin <= 24'd00025938;
                12'd0482: logsin <= 24'd00026047;
                12'd0483: logsin <= 24'd00026155;
                12'd0484: logsin <= 24'd00026264;
                12'd0485: logsin <= 24'd00026374;
                12'd0486: logsin <= 24'd00026483;
                12'd0487: logsin <= 24'd00026593;
                12'd0488: logsin <= 24'd00026702;
                12'd0489: logsin <= 24'd00026812;
                12'd0490: logsin <= 24'd00026923;
                12'd0491: logsin <= 24'd00027033;
                12'd0492: logsin <= 24'd00027144;
                12'd0493: logsin <= 24'd00027255;
                12'd0494: logsin <= 24'd00027366;
                12'd0495: logsin <= 24'd00027478;
                12'd0496: logsin <= 24'd00027590;
                12'd0497: logsin <= 24'd00027701;
                12'd0498: logsin <= 24'd00027814;
                12'd0499: logsin <= 24'd00027926;
                12'd0500: logsin <= 24'd00028039;
                12'd0501: logsin <= 24'd00028152;
                12'd0502: logsin <= 24'd00028265;
                12'd0503: logsin <= 24'd00028378;
                12'd0504: logsin <= 24'd00028491;
                12'd0505: logsin <= 24'd00028605;
                12'd0506: logsin <= 24'd00028719;
                12'd0507: logsin <= 24'd00028833;
                12'd0508: logsin <= 24'd00028948;
                12'd0509: logsin <= 24'd00029063;
                12'd0510: logsin <= 24'd00029178;
                12'd0511: logsin <= 24'd00029293;
                12'd0512: logsin <= 24'd00029408;
                12'd0513: logsin <= 24'd00029524;
                12'd0514: logsin <= 24'd00029640;
                12'd0515: logsin <= 24'd00029756;
                12'd0516: logsin <= 24'd00029872;
                12'd0517: logsin <= 24'd00029989;
                12'd0518: logsin <= 24'd00030105;
                12'd0519: logsin <= 24'd00030222;
                12'd0520: logsin <= 24'd00030340;
                12'd0521: logsin <= 24'd00030457;
                12'd0522: logsin <= 24'd00030575;
                12'd0523: logsin <= 24'd00030693;
                12'd0524: logsin <= 24'd00030811;
                12'd0525: logsin <= 24'd00030929;
                12'd0526: logsin <= 24'd00031048;
                12'd0527: logsin <= 24'd00031167;
                12'd0528: logsin <= 24'd00031286;
                12'd0529: logsin <= 24'd00031405;
                12'd0530: logsin <= 24'd00031525;
                12'd0531: logsin <= 24'd00031645;
                12'd0532: logsin <= 24'd00031765;
                12'd0533: logsin <= 24'd00031885;
                12'd0534: logsin <= 24'd00032006;
                12'd0535: logsin <= 24'd00032126;
                12'd0536: logsin <= 24'd00032247;
                12'd0537: logsin <= 24'd00032368;
                12'd0538: logsin <= 24'd00032490;
                12'd0539: logsin <= 24'd00032611;
                12'd0540: logsin <= 24'd00032733;
                12'd0541: logsin <= 24'd00032855;
                12'd0542: logsin <= 24'd00032978;
                12'd0543: logsin <= 24'd00033100;
                12'd0544: logsin <= 24'd00033223;
                12'd0545: logsin <= 24'd00033346;
                12'd0546: logsin <= 24'd00033470;
                12'd0547: logsin <= 24'd00033593;
                12'd0548: logsin <= 24'd00033717;
                12'd0549: logsin <= 24'd00033841;
                12'd0550: logsin <= 24'd00033965;
                12'd0551: logsin <= 24'd00034089;
                12'd0552: logsin <= 24'd00034214;
                12'd0553: logsin <= 24'd00034339;
                12'd0554: logsin <= 24'd00034464;
                12'd0555: logsin <= 24'd00034590;
                12'd0556: logsin <= 24'd00034715;
                12'd0557: logsin <= 24'd00034841;
                12'd0558: logsin <= 24'd00034967;
                12'd0559: logsin <= 24'd00035093;
                12'd0560: logsin <= 24'd00035220;
                12'd0561: logsin <= 24'd00035347;
                12'd0562: logsin <= 24'd00035474;
                12'd0563: logsin <= 24'd00035601;
                12'd0564: logsin <= 24'd00035728;
                12'd0565: logsin <= 24'd00035856;
                12'd0566: logsin <= 24'd00035984;
                12'd0567: logsin <= 24'd00036112;
                12'd0568: logsin <= 24'd00036241;
                12'd0569: logsin <= 24'd00036369;
                12'd0570: logsin <= 24'd00036498;
                12'd0571: logsin <= 24'd00036627;
                12'd0572: logsin <= 24'd00036757;
                12'd0573: logsin <= 24'd00036886;
                12'd0574: logsin <= 24'd00037016;
                12'd0575: logsin <= 24'd00037146;
                12'd0576: logsin <= 24'd00037276;
                12'd0577: logsin <= 24'd00037407;
                12'd0578: logsin <= 24'd00037538;
                12'd0579: logsin <= 24'd00037669;
                12'd0580: logsin <= 24'd00037800;
                12'd0581: logsin <= 24'd00037931;
                12'd0582: logsin <= 24'd00038063;
                12'd0583: logsin <= 24'd00038195;
                12'd0584: logsin <= 24'd00038327;
                12'd0585: logsin <= 24'd00038459;
                12'd0586: logsin <= 24'd00038592;
                12'd0587: logsin <= 24'd00038725;
                12'd0588: logsin <= 24'd00038858;
                12'd0589: logsin <= 24'd00038991;
                12'd0590: logsin <= 24'd00039125;
                12'd0591: logsin <= 24'd00039259;
                12'd0592: logsin <= 24'd00039393;
                12'd0593: logsin <= 24'd00039527;
                12'd0594: logsin <= 24'd00039661;
                12'd0595: logsin <= 24'd00039796;
                12'd0596: logsin <= 24'd00039931;
                12'd0597: logsin <= 24'd00040066;
                12'd0598: logsin <= 24'd00040202;
                12'd0599: logsin <= 24'd00040337;
                12'd0600: logsin <= 24'd00040473;
                12'd0601: logsin <= 24'd00040609;
                12'd0602: logsin <= 24'd00040746;
                12'd0603: logsin <= 24'd00040882;
                12'd0604: logsin <= 24'd00041019;
                12'd0605: logsin <= 24'd00041156;
                12'd0606: logsin <= 24'd00041293;
                12'd0607: logsin <= 24'd00041431;
                12'd0608: logsin <= 24'd00041569;
                12'd0609: logsin <= 24'd00041707;
                12'd0610: logsin <= 24'd00041845;
                12'd0611: logsin <= 24'd00041983;
                12'd0612: logsin <= 24'd00042122;
                12'd0613: logsin <= 24'd00042261;
                12'd0614: logsin <= 24'd00042400;
                12'd0615: logsin <= 24'd00042540;
                12'd0616: logsin <= 24'd00042679;
                12'd0617: logsin <= 24'd00042819;
                12'd0618: logsin <= 24'd00042959;
                12'd0619: logsin <= 24'd00043100;
                12'd0620: logsin <= 24'd00043240;
                12'd0621: logsin <= 24'd00043381;
                12'd0622: logsin <= 24'd00043522;
                12'd0623: logsin <= 24'd00043664;
                12'd0624: logsin <= 24'd00043805;
                12'd0625: logsin <= 24'd00043947;
                12'd0626: logsin <= 24'd00044089;
                12'd0627: logsin <= 24'd00044231;
                12'd0628: logsin <= 24'd00044374;
                12'd0629: logsin <= 24'd00044516;
                12'd0630: logsin <= 24'd00044659;
                12'd0631: logsin <= 24'd00044803;
                12'd0632: logsin <= 24'd00044946;
                12'd0633: logsin <= 24'd00045090;
                12'd0634: logsin <= 24'd00045234;
                12'd0635: logsin <= 24'd00045378;
                12'd0636: logsin <= 24'd00045522;
                12'd0637: logsin <= 24'd00045667;
                12'd0638: logsin <= 24'd00045811;
                12'd0639: logsin <= 24'd00045957;
                12'd0640: logsin <= 24'd00046102;
                12'd0641: logsin <= 24'd00046247;
                12'd0642: logsin <= 24'd00046393;
                12'd0643: logsin <= 24'd00046539;
                12'd0644: logsin <= 24'd00046686;
                12'd0645: logsin <= 24'd00046832;
                12'd0646: logsin <= 24'd00046979;
                12'd0647: logsin <= 24'd00047126;
                12'd0648: logsin <= 24'd00047273;
                12'd0649: logsin <= 24'd00047420;
                12'd0650: logsin <= 24'd00047568;
                12'd0651: logsin <= 24'd00047716;
                12'd0652: logsin <= 24'd00047864;
                12'd0653: logsin <= 24'd00048013;
                12'd0654: logsin <= 24'd00048161;
                12'd0655: logsin <= 24'd00048310;
                12'd0656: logsin <= 24'd00048459;
                12'd0657: logsin <= 24'd00048609;
                12'd0658: logsin <= 24'd00048758;
                12'd0659: logsin <= 24'd00048908;
                12'd0660: logsin <= 24'd00049058;
                12'd0661: logsin <= 24'd00049208;
                12'd0662: logsin <= 24'd00049359;
                12'd0663: logsin <= 24'd00049510;
                12'd0664: logsin <= 24'd00049661;
                12'd0665: logsin <= 24'd00049812;
                12'd0666: logsin <= 24'd00049963;
                12'd0667: logsin <= 24'd00050115;
                12'd0668: logsin <= 24'd00050267;
                12'd0669: logsin <= 24'd00050419;
                12'd0670: logsin <= 24'd00050572;
                12'd0671: logsin <= 24'd00050724;
                12'd0672: logsin <= 24'd00050877;
                12'd0673: logsin <= 24'd00051030;
                12'd0674: logsin <= 24'd00051184;
                12'd0675: logsin <= 24'd00051337;
                12'd0676: logsin <= 24'd00051491;
                12'd0677: logsin <= 24'd00051645;
                12'd0678: logsin <= 24'd00051800;
                12'd0679: logsin <= 24'd00051954;
                12'd0680: logsin <= 24'd00052109;
                12'd0681: logsin <= 24'd00052264;
                12'd0682: logsin <= 24'd00052419;
                12'd0683: logsin <= 24'd00052575;
                12'd0684: logsin <= 24'd00052731;
                12'd0685: logsin <= 24'd00052887;
                12'd0686: logsin <= 24'd00053043;
                12'd0687: logsin <= 24'd00053199;
                12'd0688: logsin <= 24'd00053356;
                12'd0689: logsin <= 24'd00053513;
                12'd0690: logsin <= 24'd00053670;
                12'd0691: logsin <= 24'd00053828;
                12'd0692: logsin <= 24'd00053985;
                12'd0693: logsin <= 24'd00054143;
                12'd0694: logsin <= 24'd00054301;
                12'd0695: logsin <= 24'd00054460;
                12'd0696: logsin <= 24'd00054618;
                12'd0697: logsin <= 24'd00054777;
                12'd0698: logsin <= 24'd00054936;
                12'd0699: logsin <= 24'd00055096;
                12'd0700: logsin <= 24'd00055255;
                12'd0701: logsin <= 24'd00055415;
                12'd0702: logsin <= 24'd00055575;
                12'd0703: logsin <= 24'd00055736;
                12'd0704: logsin <= 24'd00055896;
                12'd0705: logsin <= 24'd00056057;
                12'd0706: logsin <= 24'd00056218;
                12'd0707: logsin <= 24'd00056379;
                12'd0708: logsin <= 24'd00056541;
                12'd0709: logsin <= 24'd00056702;
                12'd0710: logsin <= 24'd00056864;
                12'd0711: logsin <= 24'd00057027;
                12'd0712: logsin <= 24'd00057189;
                12'd0713: logsin <= 24'd00057352;
                12'd0714: logsin <= 24'd00057515;
                12'd0715: logsin <= 24'd00057678;
                12'd0716: logsin <= 24'd00057841;
                12'd0717: logsin <= 24'd00058005;
                12'd0718: logsin <= 24'd00058169;
                12'd0719: logsin <= 24'd00058333;
                12'd0720: logsin <= 24'd00058497;
                12'd0721: logsin <= 24'd00058662;
                12'd0722: logsin <= 24'd00058827;
                12'd0723: logsin <= 24'd00058992;
                12'd0724: logsin <= 24'd00059157;
                12'd0725: logsin <= 24'd00059323;
                12'd0726: logsin <= 24'd00059489;
                12'd0727: logsin <= 24'd00059655;
                12'd0728: logsin <= 24'd00059821;
                12'd0729: logsin <= 24'd00059988;
                12'd0730: logsin <= 24'd00060155;
                12'd0731: logsin <= 24'd00060322;
                12'd0732: logsin <= 24'd00060489;
                12'd0733: logsin <= 24'd00060656;
                12'd0734: logsin <= 24'd00060824;
                12'd0735: logsin <= 24'd00060992;
                12'd0736: logsin <= 24'd00061160;
                12'd0737: logsin <= 24'd00061329;
                12'd0738: logsin <= 24'd00061498;
                12'd0739: logsin <= 24'd00061667;
                12'd0740: logsin <= 24'd00061836;
                12'd0741: logsin <= 24'd00062005;
                12'd0742: logsin <= 24'd00062175;
                12'd0743: logsin <= 24'd00062345;
                12'd0744: logsin <= 24'd00062515;
                12'd0745: logsin <= 24'd00062685;
                12'd0746: logsin <= 24'd00062856;
                12'd0747: logsin <= 24'd00063027;
                12'd0748: logsin <= 24'd00063198;
                12'd0749: logsin <= 24'd00063369;
                12'd0750: logsin <= 24'd00063541;
                12'd0751: logsin <= 24'd00063713;
                12'd0752: logsin <= 24'd00063885;
                12'd0753: logsin <= 24'd00064057;
                12'd0754: logsin <= 24'd00064230;
                12'd0755: logsin <= 24'd00064403;
                12'd0756: logsin <= 24'd00064576;
                12'd0757: logsin <= 24'd00064749;
                12'd0758: logsin <= 24'd00064923;
                12'd0759: logsin <= 24'd00065097;
                12'd0760: logsin <= 24'd00065271;
                12'd0761: logsin <= 24'd00065445;
                12'd0762: logsin <= 24'd00065619;
                12'd0763: logsin <= 24'd00065794;
                12'd0764: logsin <= 24'd00065969;
                12'd0765: logsin <= 24'd00066144;
                12'd0766: logsin <= 24'd00066320;
                12'd0767: logsin <= 24'd00066496;
                12'd0768: logsin <= 24'd00066672;
                12'd0769: logsin <= 24'd00066848;
                12'd0770: logsin <= 24'd00067024;
                12'd0771: logsin <= 24'd00067201;
                12'd0772: logsin <= 24'd00067378;
                12'd0773: logsin <= 24'd00067555;
                12'd0774: logsin <= 24'd00067733;
                12'd0775: logsin <= 24'd00067910;
                12'd0776: logsin <= 24'd00068088;
                12'd0777: logsin <= 24'd00068266;
                12'd0778: logsin <= 24'd00068445;
                12'd0779: logsin <= 24'd00068624;
                12'd0780: logsin <= 24'd00068802;
                12'd0781: logsin <= 24'd00068982;
                12'd0782: logsin <= 24'd00069161;
                12'd0783: logsin <= 24'd00069341;
                12'd0784: logsin <= 24'd00069521;
                12'd0785: logsin <= 24'd00069701;
                12'd0786: logsin <= 24'd00069881;
                12'd0787: logsin <= 24'd00070062;
                12'd0788: logsin <= 24'd00070242;
                12'd0789: logsin <= 24'd00070424;
                12'd0790: logsin <= 24'd00070605;
                12'd0791: logsin <= 24'd00070786;
                12'd0792: logsin <= 24'd00070968;
                12'd0793: logsin <= 24'd00071150;
                12'd0794: logsin <= 24'd00071333;
                12'd0795: logsin <= 24'd00071515;
                12'd0796: logsin <= 24'd00071698;
                12'd0797: logsin <= 24'd00071881;
                12'd0798: logsin <= 24'd00072064;
                12'd0799: logsin <= 24'd00072248;
                12'd0800: logsin <= 24'd00072432;
                12'd0801: logsin <= 24'd00072616;
                12'd0802: logsin <= 24'd00072800;
                12'd0803: logsin <= 24'd00072985;
                12'd0804: logsin <= 24'd00073169;
                12'd0805: logsin <= 24'd00073354;
                12'd0806: logsin <= 24'd00073540;
                12'd0807: logsin <= 24'd00073725;
                12'd0808: logsin <= 24'd00073911;
                12'd0809: logsin <= 24'd00074097;
                12'd0810: logsin <= 24'd00074283;
                12'd0811: logsin <= 24'd00074470;
                12'd0812: logsin <= 24'd00074656;
                12'd0813: logsin <= 24'd00074843;
                12'd0814: logsin <= 24'd00075031;
                12'd0815: logsin <= 24'd00075218;
                12'd0816: logsin <= 24'd00075406;
                12'd0817: logsin <= 24'd00075594;
                12'd0818: logsin <= 24'd00075782;
                12'd0819: logsin <= 24'd00075970;
                12'd0820: logsin <= 24'd00076159;
                12'd0821: logsin <= 24'd00076348;
                12'd0822: logsin <= 24'd00076537;
                12'd0823: logsin <= 24'd00076727;
                12'd0824: logsin <= 24'd00076916;
                12'd0825: logsin <= 24'd00077106;
                12'd0826: logsin <= 24'd00077296;
                12'd0827: logsin <= 24'd00077487;
                12'd0828: logsin <= 24'd00077677;
                12'd0829: logsin <= 24'd00077868;
                12'd0830: logsin <= 24'd00078060;
                12'd0831: logsin <= 24'd00078251;
                12'd0832: logsin <= 24'd00078443;
                12'd0833: logsin <= 24'd00078635;
                12'd0834: logsin <= 24'd00078827;
                12'd0835: logsin <= 24'd00079019;
                12'd0836: logsin <= 24'd00079212;
                12'd0837: logsin <= 24'd00079405;
                12'd0838: logsin <= 24'd00079598;
                12'd0839: logsin <= 24'd00079791;
                12'd0840: logsin <= 24'd00079985;
                12'd0841: logsin <= 24'd00080179;
                12'd0842: logsin <= 24'd00080373;
                12'd0843: logsin <= 24'd00080567;
                12'd0844: logsin <= 24'd00080762;
                12'd0845: logsin <= 24'd00080957;
                12'd0846: logsin <= 24'd00081152;
                12'd0847: logsin <= 24'd00081347;
                12'd0848: logsin <= 24'd00081543;
                12'd0849: logsin <= 24'd00081739;
                12'd0850: logsin <= 24'd00081935;
                12'd0851: logsin <= 24'd00082131;
                12'd0852: logsin <= 24'd00082328;
                12'd0853: logsin <= 24'd00082524;
                12'd0854: logsin <= 24'd00082722;
                12'd0855: logsin <= 24'd00082919;
                12'd0856: logsin <= 24'd00083116;
                12'd0857: logsin <= 24'd00083314;
                12'd0858: logsin <= 24'd00083512;
                12'd0859: logsin <= 24'd00083711;
                12'd0860: logsin <= 24'd00083909;
                12'd0861: logsin <= 24'd00084108;
                12'd0862: logsin <= 24'd00084307;
                12'd0863: logsin <= 24'd00084507;
                12'd0864: logsin <= 24'd00084706;
                12'd0865: logsin <= 24'd00084906;
                12'd0866: logsin <= 24'd00085106;
                12'd0867: logsin <= 24'd00085306;
                12'd0868: logsin <= 24'd00085507;
                12'd0869: logsin <= 24'd00085708;
                12'd0870: logsin <= 24'd00085909;
                12'd0871: logsin <= 24'd00086110;
                12'd0872: logsin <= 24'd00086312;
                12'd0873: logsin <= 24'd00086514;
                12'd0874: logsin <= 24'd00086716;
                12'd0875: logsin <= 24'd00086918;
                12'd0876: logsin <= 24'd00087121;
                12'd0877: logsin <= 24'd00087323;
                12'd0878: logsin <= 24'd00087526;
                12'd0879: logsin <= 24'd00087730;
                12'd0880: logsin <= 24'd00087933;
                12'd0881: logsin <= 24'd00088137;
                12'd0882: logsin <= 24'd00088341;
                12'd0883: logsin <= 24'd00088546;
                12'd0884: logsin <= 24'd00088750;
                12'd0885: logsin <= 24'd00088955;
                12'd0886: logsin <= 24'd00089160;
                12'd0887: logsin <= 24'd00089365;
                12'd0888: logsin <= 24'd00089571;
                12'd0889: logsin <= 24'd00089777;
                12'd0890: logsin <= 24'd00089983;
                12'd0891: logsin <= 24'd00090189;
                12'd0892: logsin <= 24'd00090396;
                12'd0893: logsin <= 24'd00090603;
                12'd0894: logsin <= 24'd00090810;
                12'd0895: logsin <= 24'd00091017;
                12'd0896: logsin <= 24'd00091225;
                12'd0897: logsin <= 24'd00091432;
                12'd0898: logsin <= 24'd00091640;
                12'd0899: logsin <= 24'd00091849;
                12'd0900: logsin <= 24'd00092057;
                12'd0901: logsin <= 24'd00092266;
                12'd0902: logsin <= 24'd00092475;
                12'd0903: logsin <= 24'd00092685;
                12'd0904: logsin <= 24'd00092894;
                12'd0905: logsin <= 24'd00093104;
                12'd0906: logsin <= 24'd00093314;
                12'd0907: logsin <= 24'd00093524;
                12'd0908: logsin <= 24'd00093735;
                12'd0909: logsin <= 24'd00093946;
                12'd0910: logsin <= 24'd00094157;
                12'd0911: logsin <= 24'd00094368;
                12'd0912: logsin <= 24'd00094580;
                12'd0913: logsin <= 24'd00094792;
                12'd0914: logsin <= 24'd00095004;
                12'd0915: logsin <= 24'd00095216;
                12'd0916: logsin <= 24'd00095429;
                12'd0917: logsin <= 24'd00095642;
                12'd0918: logsin <= 24'd00095855;
                12'd0919: logsin <= 24'd00096068;
                12'd0920: logsin <= 24'd00096282;
                12'd0921: logsin <= 24'd00096496;
                12'd0922: logsin <= 24'd00096710;
                12'd0923: logsin <= 24'd00096924;
                12'd0924: logsin <= 24'd00097139;
                12'd0925: logsin <= 24'd00097354;
                12'd0926: logsin <= 24'd00097569;
                12'd0927: logsin <= 24'd00097784;
                12'd0928: logsin <= 24'd00098000;
                12'd0929: logsin <= 24'd00098216;
                12'd0930: logsin <= 24'd00098432;
                12'd0931: logsin <= 24'd00098648;
                12'd0932: logsin <= 24'd00098865;
                12'd0933: logsin <= 24'd00099082;
                12'd0934: logsin <= 24'd00099299;
                12'd0935: logsin <= 24'd00099517;
                12'd0936: logsin <= 24'd00099734;
                12'd0937: logsin <= 24'd00099952;
                12'd0938: logsin <= 24'd00100170;
                12'd0939: logsin <= 24'd00100389;
                12'd0940: logsin <= 24'd00100607;
                12'd0941: logsin <= 24'd00100826;
                12'd0942: logsin <= 24'd00101046;
                12'd0943: logsin <= 24'd00101265;
                12'd0944: logsin <= 24'd00101485;
                12'd0945: logsin <= 24'd00101705;
                12'd0946: logsin <= 24'd00101925;
                12'd0947: logsin <= 24'd00102145;
                12'd0948: logsin <= 24'd00102366;
                12'd0949: logsin <= 24'd00102587;
                12'd0950: logsin <= 24'd00102808;
                12'd0951: logsin <= 24'd00103030;
                12'd0952: logsin <= 24'd00103252;
                12'd0953: logsin <= 24'd00103474;
                12'd0954: logsin <= 24'd00103696;
                12'd0955: logsin <= 24'd00103918;
                12'd0956: logsin <= 24'd00104141;
                12'd0957: logsin <= 24'd00104364;
                12'd0958: logsin <= 24'd00104587;
                12'd0959: logsin <= 24'd00104811;
                12'd0960: logsin <= 24'd00105035;
                12'd0961: logsin <= 24'd00105259;
                12'd0962: logsin <= 24'd00105483;
                12'd0963: logsin <= 24'd00105708;
                12'd0964: logsin <= 24'd00105932;
                12'd0965: logsin <= 24'd00106157;
                12'd0966: logsin <= 24'd00106383;
                12'd0967: logsin <= 24'd00106608;
                12'd0968: logsin <= 24'd00106834;
                12'd0969: logsin <= 24'd00107060;
                12'd0970: logsin <= 24'd00107287;
                12'd0971: logsin <= 24'd00107513;
                12'd0972: logsin <= 24'd00107740;
                12'd0973: logsin <= 24'd00107967;
                12'd0974: logsin <= 24'd00108195;
                12'd0975: logsin <= 24'd00108422;
                12'd0976: logsin <= 24'd00108650;
                12'd0977: logsin <= 24'd00108878;
                12'd0978: logsin <= 24'd00109107;
                12'd0979: logsin <= 24'd00109335;
                12'd0980: logsin <= 24'd00109564;
                12'd0981: logsin <= 24'd00109793;
                12'd0982: logsin <= 24'd00110023;
                12'd0983: logsin <= 24'd00110252;
                12'd0984: logsin <= 24'd00110482;
                12'd0985: logsin <= 24'd00110713;
                12'd0986: logsin <= 24'd00110943;
                12'd0987: logsin <= 24'd00111174;
                12'd0988: logsin <= 24'd00111405;
                12'd0989: logsin <= 24'd00111636;
                12'd0990: logsin <= 24'd00111867;
                12'd0991: logsin <= 24'd00112099;
                12'd0992: logsin <= 24'd00112331;
                12'd0993: logsin <= 24'd00112563;
                12'd0994: logsin <= 24'd00112796;
                12'd0995: logsin <= 24'd00113029;
                12'd0996: logsin <= 24'd00113262;
                12'd0997: logsin <= 24'd00113495;
                12'd0998: logsin <= 24'd00113729;
                12'd0999: logsin <= 24'd00113962;
                12'd1000: logsin <= 24'd00114197;
                12'd1001: logsin <= 24'd00114431;
                12'd1002: logsin <= 24'd00114665;
                12'd1003: logsin <= 24'd00114900;
                12'd1004: logsin <= 24'd00115135;
                12'd1005: logsin <= 24'd00115371;
                12'd1006: logsin <= 24'd00115606;
                12'd1007: logsin <= 24'd00115842;
                12'd1008: logsin <= 24'd00116078;
                12'd1009: logsin <= 24'd00116315;
                12'd1010: logsin <= 24'd00116551;
                12'd1011: logsin <= 24'd00116788;
                12'd1012: logsin <= 24'd00117026;
                12'd1013: logsin <= 24'd00117263;
                12'd1014: logsin <= 24'd00117501;
                12'd1015: logsin <= 24'd00117739;
                12'd1016: logsin <= 24'd00117977;
                12'd1017: logsin <= 24'd00118215;
                12'd1018: logsin <= 24'd00118454;
                12'd1019: logsin <= 24'd00118693;
                12'd1020: logsin <= 24'd00118932;
                12'd1021: logsin <= 24'd00119172;
                12'd1022: logsin <= 24'd00119412;
                12'd1023: logsin <= 24'd00119652;
                12'd1024: logsin <= 24'd00119892;
                12'd1025: logsin <= 24'd00120133;
                12'd1026: logsin <= 24'd00120373;
                12'd1027: logsin <= 24'd00120615;
                12'd1028: logsin <= 24'd00120856;
                12'd1029: logsin <= 24'd00121097;
                12'd1030: logsin <= 24'd00121339;
                12'd1031: logsin <= 24'd00121581;
                12'd1032: logsin <= 24'd00121824;
                12'd1033: logsin <= 24'd00122067;
                12'd1034: logsin <= 24'd00122309;
                12'd1035: logsin <= 24'd00122553;
                12'd1036: logsin <= 24'd00122796;
                12'd1037: logsin <= 24'd00123040;
                12'd1038: logsin <= 24'd00123284;
                12'd1039: logsin <= 24'd00123528;
                12'd1040: logsin <= 24'd00123772;
                12'd1041: logsin <= 24'd00124017;
                12'd1042: logsin <= 24'd00124262;
                12'd1043: logsin <= 24'd00124507;
                12'd1044: logsin <= 24'd00124753;
                12'd1045: logsin <= 24'd00124999;
                12'd1046: logsin <= 24'd00125245;
                12'd1047: logsin <= 24'd00125491;
                12'd1048: logsin <= 24'd00125738;
                12'd1049: logsin <= 24'd00125985;
                12'd1050: logsin <= 24'd00126232;
                12'd1051: logsin <= 24'd00126479;
                12'd1052: logsin <= 24'd00126727;
                12'd1053: logsin <= 24'd00126975;
                12'd1054: logsin <= 24'd00127223;
                12'd1055: logsin <= 24'd00127471;
                12'd1056: logsin <= 24'd00127720;
                12'd1057: logsin <= 24'd00127969;
                12'd1058: logsin <= 24'd00128218;
                12'd1059: logsin <= 24'd00128467;
                12'd1060: logsin <= 24'd00128717;
                12'd1061: logsin <= 24'd00128967;
                12'd1062: logsin <= 24'd00129217;
                12'd1063: logsin <= 24'd00129468;
                12'd1064: logsin <= 24'd00129719;
                12'd1065: logsin <= 24'd00129970;
                12'd1066: logsin <= 24'd00130221;
                12'd1067: logsin <= 24'd00130473;
                12'd1068: logsin <= 24'd00130725;
                12'd1069: logsin <= 24'd00130977;
                12'd1070: logsin <= 24'd00131229;
                12'd1071: logsin <= 24'd00131482;
                12'd1072: logsin <= 24'd00131735;
                12'd1073: logsin <= 24'd00131988;
                12'd1074: logsin <= 24'd00132241;
                12'd1075: logsin <= 24'd00132495;
                12'd1076: logsin <= 24'd00132749;
                12'd1077: logsin <= 24'd00133003;
                12'd1078: logsin <= 24'd00133258;
                12'd1079: logsin <= 24'd00133513;
                12'd1080: logsin <= 24'd00133768;
                12'd1081: logsin <= 24'd00134023;
                12'd1082: logsin <= 24'd00134278;
                12'd1083: logsin <= 24'd00134534;
                12'd1084: logsin <= 24'd00134790;
                12'd1085: logsin <= 24'd00135047;
                12'd1086: logsin <= 24'd00135303;
                12'd1087: logsin <= 24'd00135560;
                12'd1088: logsin <= 24'd00135817;
                12'd1089: logsin <= 24'd00136075;
                12'd1090: logsin <= 24'd00136332;
                12'd1091: logsin <= 24'd00136590;
                12'd1092: logsin <= 24'd00136849;
                12'd1093: logsin <= 24'd00137107;
                12'd1094: logsin <= 24'd00137366;
                12'd1095: logsin <= 24'd00137625;
                12'd1096: logsin <= 24'd00137884;
                12'd1097: logsin <= 24'd00138144;
                12'd1098: logsin <= 24'd00138404;
                12'd1099: logsin <= 24'd00138664;
                12'd1100: logsin <= 24'd00138924;
                12'd1101: logsin <= 24'd00139185;
                12'd1102: logsin <= 24'd00139446;
                12'd1103: logsin <= 24'd00139707;
                12'd1104: logsin <= 24'd00139968;
                12'd1105: logsin <= 24'd00140230;
                12'd1106: logsin <= 24'd00140492;
                12'd1107: logsin <= 24'd00140754;
                12'd1108: logsin <= 24'd00141017;
                12'd1109: logsin <= 24'd00141279;
                12'd1110: logsin <= 24'd00141542;
                12'd1111: logsin <= 24'd00141806;
                12'd1112: logsin <= 24'd00142069;
                12'd1113: logsin <= 24'd00142333;
                12'd1114: logsin <= 24'd00142597;
                12'd1115: logsin <= 24'd00142862;
                12'd1116: logsin <= 24'd00143126;
                12'd1117: logsin <= 24'd00143391;
                12'd1118: logsin <= 24'd00143656;
                12'd1119: logsin <= 24'd00143922;
                12'd1120: logsin <= 24'd00144188;
                12'd1121: logsin <= 24'd00144454;
                12'd1122: logsin <= 24'd00144720;
                12'd1123: logsin <= 24'd00144986;
                12'd1124: logsin <= 24'd00145253;
                12'd1125: logsin <= 24'd00145520;
                12'd1126: logsin <= 24'd00145788;
                12'd1127: logsin <= 24'd00146055;
                12'd1128: logsin <= 24'd00146323;
                12'd1129: logsin <= 24'd00146591;
                12'd1130: logsin <= 24'd00146860;
                12'd1131: logsin <= 24'd00147128;
                12'd1132: logsin <= 24'd00147397;
                12'd1133: logsin <= 24'd00147666;
                12'd1134: logsin <= 24'd00147936;
                12'd1135: logsin <= 24'd00148206;
                12'd1136: logsin <= 24'd00148476;
                12'd1137: logsin <= 24'd00148746;
                12'd1138: logsin <= 24'd00149017;
                12'd1139: logsin <= 24'd00149288;
                12'd1140: logsin <= 24'd00149559;
                12'd1141: logsin <= 24'd00149830;
                12'd1142: logsin <= 24'd00150102;
                12'd1143: logsin <= 24'd00150374;
                12'd1144: logsin <= 24'd00150646;
                12'd1145: logsin <= 24'd00150918;
                12'd1146: logsin <= 24'd00151191;
                12'd1147: logsin <= 24'd00151464;
                12'd1148: logsin <= 24'd00151737;
                12'd1149: logsin <= 24'd00152011;
                12'd1150: logsin <= 24'd00152285;
                12'd1151: logsin <= 24'd00152559;
                12'd1152: logsin <= 24'd00152833;
                12'd1153: logsin <= 24'd00153108;
                12'd1154: logsin <= 24'd00153383;
                12'd1155: logsin <= 24'd00153658;
                12'd1156: logsin <= 24'd00153934;
                12'd1157: logsin <= 24'd00154209;
                12'd1158: logsin <= 24'd00154485;
                12'd1159: logsin <= 24'd00154762;
                12'd1160: logsin <= 24'd00155038;
                12'd1161: logsin <= 24'd00155315;
                12'd1162: logsin <= 24'd00155592;
                12'd1163: logsin <= 24'd00155870;
                12'd1164: logsin <= 24'd00156147;
                12'd1165: logsin <= 24'd00156425;
                12'd1166: logsin <= 24'd00156703;
                12'd1167: logsin <= 24'd00156982;
                12'd1168: logsin <= 24'd00157261;
                12'd1169: logsin <= 24'd00157540;
                12'd1170: logsin <= 24'd00157819;
                12'd1171: logsin <= 24'd00158099;
                12'd1172: logsin <= 24'd00158378;
                12'd1173: logsin <= 24'd00158659;
                12'd1174: logsin <= 24'd00158939;
                12'd1175: logsin <= 24'd00159220;
                12'd1176: logsin <= 24'd00159501;
                12'd1177: logsin <= 24'd00159782;
                12'd1178: logsin <= 24'd00160063;
                12'd1179: logsin <= 24'd00160345;
                12'd1180: logsin <= 24'd00160627;
                12'd1181: logsin <= 24'd00160909;
                12'd1182: logsin <= 24'd00161192;
                12'd1183: logsin <= 24'd00161475;
                12'd1184: logsin <= 24'd00161758;
                12'd1185: logsin <= 24'd00162042;
                12'd1186: logsin <= 24'd00162325;
                12'd1187: logsin <= 24'd00162609;
                12'd1188: logsin <= 24'd00162893;
                12'd1189: logsin <= 24'd00163178;
                12'd1190: logsin <= 24'd00163463;
                12'd1191: logsin <= 24'd00163748;
                12'd1192: logsin <= 24'd00164033;
                12'd1193: logsin <= 24'd00164319;
                12'd1194: logsin <= 24'd00164605;
                12'd1195: logsin <= 24'd00164891;
                12'd1196: logsin <= 24'd00165177;
                12'd1197: logsin <= 24'd00165464;
                12'd1198: logsin <= 24'd00165751;
                12'd1199: logsin <= 24'd00166038;
                12'd1200: logsin <= 24'd00166326;
                12'd1201: logsin <= 24'd00166614;
                12'd1202: logsin <= 24'd00166902;
                12'd1203: logsin <= 24'd00167190;
                12'd1204: logsin <= 24'd00167479;
                12'd1205: logsin <= 24'd00167768;
                12'd1206: logsin <= 24'd00168057;
                12'd1207: logsin <= 24'd00168347;
                12'd1208: logsin <= 24'd00168637;
                12'd1209: logsin <= 24'd00168927;
                12'd1210: logsin <= 24'd00169217;
                12'd1211: logsin <= 24'd00169508;
                12'd1212: logsin <= 24'd00169799;
                12'd1213: logsin <= 24'd00170090;
                12'd1214: logsin <= 24'd00170381;
                12'd1215: logsin <= 24'd00170673;
                12'd1216: logsin <= 24'd00170965;
                12'd1217: logsin <= 24'd00171257;
                12'd1218: logsin <= 24'd00171550;
                12'd1219: logsin <= 24'd00171843;
                12'd1220: logsin <= 24'd00172136;
                12'd1221: logsin <= 24'd00172429;
                12'd1222: logsin <= 24'd00172723;
                12'd1223: logsin <= 24'd00173017;
                12'd1224: logsin <= 24'd00173311;
                12'd1225: logsin <= 24'd00173606;
                12'd1226: logsin <= 24'd00173900;
                12'd1227: logsin <= 24'd00174196;
                12'd1228: logsin <= 24'd00174491;
                12'd1229: logsin <= 24'd00174787;
                12'd1230: logsin <= 24'd00175083;
                12'd1231: logsin <= 24'd00175379;
                12'd1232: logsin <= 24'd00175675;
                12'd1233: logsin <= 24'd00175972;
                12'd1234: logsin <= 24'd00176269;
                12'd1235: logsin <= 24'd00176566;
                12'd1236: logsin <= 24'd00176864;
                12'd1237: logsin <= 24'd00177162;
                12'd1238: logsin <= 24'd00177460;
                12'd1239: logsin <= 24'd00177759;
                12'd1240: logsin <= 24'd00178057;
                12'd1241: logsin <= 24'd00178356;
                12'd1242: logsin <= 24'd00178656;
                12'd1243: logsin <= 24'd00178955;
                12'd1244: logsin <= 24'd00179255;
                12'd1245: logsin <= 24'd00179555;
                12'd1246: logsin <= 24'd00179856;
                12'd1247: logsin <= 24'd00180156;
                12'd1248: logsin <= 24'd00180457;
                12'd1249: logsin <= 24'd00180759;
                12'd1250: logsin <= 24'd00181060;
                12'd1251: logsin <= 24'd00181362;
                12'd1252: logsin <= 24'd00181664;
                12'd1253: logsin <= 24'd00181967;
                12'd1254: logsin <= 24'd00182269;
                12'd1255: logsin <= 24'd00182572;
                12'd1256: logsin <= 24'd00182876;
                12'd1257: logsin <= 24'd00183179;
                12'd1258: logsin <= 24'd00183483;
                12'd1259: logsin <= 24'd00183787;
                12'd1260: logsin <= 24'd00184091;
                12'd1261: logsin <= 24'd00184396;
                12'd1262: logsin <= 24'd00184701;
                12'd1263: logsin <= 24'd00185006;
                12'd1264: logsin <= 24'd00185312;
                12'd1265: logsin <= 24'd00185618;
                12'd1266: logsin <= 24'd00185924;
                12'd1267: logsin <= 24'd00186230;
                12'd1268: logsin <= 24'd00186537;
                12'd1269: logsin <= 24'd00186844;
                12'd1270: logsin <= 24'd00187151;
                12'd1271: logsin <= 24'd00187459;
                12'd1272: logsin <= 24'd00187766;
                12'd1273: logsin <= 24'd00188074;
                12'd1274: logsin <= 24'd00188383;
                12'd1275: logsin <= 24'd00188691;
                12'd1276: logsin <= 24'd00189000;
                12'd1277: logsin <= 24'd00189310;
                12'd1278: logsin <= 24'd00189619;
                12'd1279: logsin <= 24'd00189929;
                12'd1280: logsin <= 24'd00190239;
                12'd1281: logsin <= 24'd00190549;
                12'd1282: logsin <= 24'd00190860;
                12'd1283: logsin <= 24'd00191171;
                12'd1284: logsin <= 24'd00191482;
                12'd1285: logsin <= 24'd00191794;
                12'd1286: logsin <= 24'd00192106;
                12'd1287: logsin <= 24'd00192418;
                12'd1288: logsin <= 24'd00192730;
                12'd1289: logsin <= 24'd00193043;
                12'd1290: logsin <= 24'd00193356;
                12'd1291: logsin <= 24'd00193669;
                12'd1292: logsin <= 24'd00193983;
                12'd1293: logsin <= 24'd00194296;
                12'd1294: logsin <= 24'd00194610;
                12'd1295: logsin <= 24'd00194925;
                12'd1296: logsin <= 24'd00195240;
                12'd1297: logsin <= 24'd00195555;
                12'd1298: logsin <= 24'd00195870;
                12'd1299: logsin <= 24'd00196185;
                12'd1300: logsin <= 24'd00196501;
                12'd1301: logsin <= 24'd00196817;
                12'd1302: logsin <= 24'd00197134;
                12'd1303: logsin <= 24'd00197450;
                12'd1304: logsin <= 24'd00197767;
                12'd1305: logsin <= 24'd00198085;
                12'd1306: logsin <= 24'd00198402;
                12'd1307: logsin <= 24'd00198720;
                12'd1308: logsin <= 24'd00199038;
                12'd1309: logsin <= 24'd00199357;
                12'd1310: logsin <= 24'd00199675;
                12'd1311: logsin <= 24'd00199994;
                12'd1312: logsin <= 24'd00200314;
                12'd1313: logsin <= 24'd00200633;
                12'd1314: logsin <= 24'd00200953;
                12'd1315: logsin <= 24'd00201273;
                12'd1316: logsin <= 24'd00201594;
                12'd1317: logsin <= 24'd00201915;
                12'd1318: logsin <= 24'd00202236;
                12'd1319: logsin <= 24'd00202557;
                12'd1320: logsin <= 24'd00202879;
                12'd1321: logsin <= 24'd00203201;
                12'd1322: logsin <= 24'd00203523;
                12'd1323: logsin <= 24'd00203845;
                12'd1324: logsin <= 24'd00204168;
                12'd1325: logsin <= 24'd00204491;
                12'd1326: logsin <= 24'd00204815;
                12'd1327: logsin <= 24'd00205138;
                12'd1328: logsin <= 24'd00205462;
                12'd1329: logsin <= 24'd00205786;
                12'd1330: logsin <= 24'd00206111;
                12'd1331: logsin <= 24'd00206436;
                12'd1332: logsin <= 24'd00206761;
                12'd1333: logsin <= 24'd00207086;
                12'd1334: logsin <= 24'd00207412;
                12'd1335: logsin <= 24'd00207738;
                12'd1336: logsin <= 24'd00208064;
                12'd1337: logsin <= 24'd00208391;
                12'd1338: logsin <= 24'd00208718;
                12'd1339: logsin <= 24'd00209045;
                12'd1340: logsin <= 24'd00209373;
                12'd1341: logsin <= 24'd00209700;
                12'd1342: logsin <= 24'd00210028;
                12'd1343: logsin <= 24'd00210357;
                12'd1344: logsin <= 24'd00210685;
                12'd1345: logsin <= 24'd00211014;
                12'd1346: logsin <= 24'd00211344;
                12'd1347: logsin <= 24'd00211673;
                12'd1348: logsin <= 24'd00212003;
                12'd1349: logsin <= 24'd00212333;
                12'd1350: logsin <= 24'd00212663;
                12'd1351: logsin <= 24'd00212994;
                12'd1352: logsin <= 24'd00213325;
                12'd1353: logsin <= 24'd00213656;
                12'd1354: logsin <= 24'd00213988;
                12'd1355: logsin <= 24'd00214320;
                12'd1356: logsin <= 24'd00214652;
                12'd1357: logsin <= 24'd00214985;
                12'd1358: logsin <= 24'd00215317;
                12'd1359: logsin <= 24'd00215650;
                12'd1360: logsin <= 24'd00215984;
                12'd1361: logsin <= 24'd00216317;
                12'd1362: logsin <= 24'd00216651;
                12'd1363: logsin <= 24'd00216986;
                12'd1364: logsin <= 24'd00217320;
                12'd1365: logsin <= 24'd00217655;
                12'd1366: logsin <= 24'd00217990;
                12'd1367: logsin <= 24'd00218326;
                12'd1368: logsin <= 24'd00218661;
                12'd1369: logsin <= 24'd00218997;
                12'd1370: logsin <= 24'd00219334;
                12'd1371: logsin <= 24'd00219670;
                12'd1372: logsin <= 24'd00220007;
                12'd1373: logsin <= 24'd00220344;
                12'd1374: logsin <= 24'd00220682;
                12'd1375: logsin <= 24'd00221020;
                12'd1376: logsin <= 24'd00221358;
                12'd1377: logsin <= 24'd00221696;
                12'd1378: logsin <= 24'd00222035;
                12'd1379: logsin <= 24'd00222374;
                12'd1380: logsin <= 24'd00222713;
                12'd1381: logsin <= 24'd00223053;
                12'd1382: logsin <= 24'd00223393;
                12'd1383: logsin <= 24'd00223733;
                12'd1384: logsin <= 24'd00224074;
                12'd1385: logsin <= 24'd00224414;
                12'd1386: logsin <= 24'd00224756;
                12'd1387: logsin <= 24'd00225097;
                12'd1388: logsin <= 24'd00225439;
                12'd1389: logsin <= 24'd00225781;
                12'd1390: logsin <= 24'd00226123;
                12'd1391: logsin <= 24'd00226466;
                12'd1392: logsin <= 24'd00226808;
                12'd1393: logsin <= 24'd00227152;
                12'd1394: logsin <= 24'd00227495;
                12'd1395: logsin <= 24'd00227839;
                12'd1396: logsin <= 24'd00228183;
                12'd1397: logsin <= 24'd00228527;
                12'd1398: logsin <= 24'd00228872;
                12'd1399: logsin <= 24'd00229217;
                12'd1400: logsin <= 24'd00229562;
                12'd1401: logsin <= 24'd00229908;
                12'd1402: logsin <= 24'd00230254;
                12'd1403: logsin <= 24'd00230600;
                12'd1404: logsin <= 24'd00230947;
                12'd1405: logsin <= 24'd00231294;
                12'd1406: logsin <= 24'd00231641;
                12'd1407: logsin <= 24'd00231988;
                12'd1408: logsin <= 24'd00232336;
                12'd1409: logsin <= 24'd00232684;
                12'd1410: logsin <= 24'd00233032;
                12'd1411: logsin <= 24'd00233381;
                12'd1412: logsin <= 24'd00233730;
                12'd1413: logsin <= 24'd00234079;
                12'd1414: logsin <= 24'd00234429;
                12'd1415: logsin <= 24'd00234778;
                12'd1416: logsin <= 24'd00235129;
                12'd1417: logsin <= 24'd00235479;
                12'd1418: logsin <= 24'd00235830;
                12'd1419: logsin <= 24'd00236181;
                12'd1420: logsin <= 24'd00236532;
                12'd1421: logsin <= 24'd00236884;
                12'd1422: logsin <= 24'd00237236;
                12'd1423: logsin <= 24'd00237588;
                12'd1424: logsin <= 24'd00237941;
                12'd1425: logsin <= 24'd00238294;
                12'd1426: logsin <= 24'd00238647;
                12'd1427: logsin <= 24'd00239000;
                12'd1428: logsin <= 24'd00239354;
                12'd1429: logsin <= 24'd00239708;
                12'd1430: logsin <= 24'd00240063;
                12'd1431: logsin <= 24'd00240417;
                12'd1432: logsin <= 24'd00240772;
                12'd1433: logsin <= 24'd00241128;
                12'd1434: logsin <= 24'd00241483;
                12'd1435: logsin <= 24'd00241839;
                12'd1436: logsin <= 24'd00242195;
                12'd1437: logsin <= 24'd00242552;
                12'd1438: logsin <= 24'd00242909;
                12'd1439: logsin <= 24'd00243266;
                12'd1440: logsin <= 24'd00243623;
                12'd1441: logsin <= 24'd00243981;
                12'd1442: logsin <= 24'd00244339;
                12'd1443: logsin <= 24'd00244698;
                12'd1444: logsin <= 24'd00245056;
                12'd1445: logsin <= 24'd00245415;
                12'd1446: logsin <= 24'd00245775;
                12'd1447: logsin <= 24'd00246134;
                12'd1448: logsin <= 24'd00246494;
                12'd1449: logsin <= 24'd00246855;
                12'd1450: logsin <= 24'd00247215;
                12'd1451: logsin <= 24'd00247576;
                12'd1452: logsin <= 24'd00247937;
                12'd1453: logsin <= 24'd00248299;
                12'd1454: logsin <= 24'd00248660;
                12'd1455: logsin <= 24'd00249022;
                12'd1456: logsin <= 24'd00249385;
                12'd1457: logsin <= 24'd00249748;
                12'd1458: logsin <= 24'd00250111;
                12'd1459: logsin <= 24'd00250474;
                12'd1460: logsin <= 24'd00250838;
                12'd1461: logsin <= 24'd00251202;
                12'd1462: logsin <= 24'd00251566;
                12'd1463: logsin <= 24'd00251930;
                12'd1464: logsin <= 24'd00252295;
                12'd1465: logsin <= 24'd00252660;
                12'd1466: logsin <= 24'd00253026;
                12'd1467: logsin <= 24'd00253392;
                12'd1468: logsin <= 24'd00253758;
                12'd1469: logsin <= 24'd00254124;
                12'd1470: logsin <= 24'd00254491;
                12'd1471: logsin <= 24'd00254858;
                12'd1472: logsin <= 24'd00255225;
                12'd1473: logsin <= 24'd00255593;
                12'd1474: logsin <= 24'd00255961;
                12'd1475: logsin <= 24'd00256329;
                12'd1476: logsin <= 24'd00256698;
                12'd1477: logsin <= 24'd00257067;
                12'd1478: logsin <= 24'd00257436;
                12'd1479: logsin <= 24'd00257806;
                12'd1480: logsin <= 24'd00258176;
                12'd1481: logsin <= 24'd00258546;
                12'd1482: logsin <= 24'd00258916;
                12'd1483: logsin <= 24'd00259287;
                12'd1484: logsin <= 24'd00259658;
                12'd1485: logsin <= 24'd00260030;
                12'd1486: logsin <= 24'd00260401;
                12'd1487: logsin <= 24'd00260774;
                12'd1488: logsin <= 24'd00261146;
                12'd1489: logsin <= 24'd00261519;
                12'd1490: logsin <= 24'd00261892;
                12'd1491: logsin <= 24'd00262265;
                12'd1492: logsin <= 24'd00262639;
                12'd1493: logsin <= 24'd00263013;
                12'd1494: logsin <= 24'd00263387;
                12'd1495: logsin <= 24'd00263761;
                12'd1496: logsin <= 24'd00264136;
                12'd1497: logsin <= 24'd00264511;
                12'd1498: logsin <= 24'd00264887;
                12'd1499: logsin <= 24'd00265263;
                12'd1500: logsin <= 24'd00265639;
                12'd1501: logsin <= 24'd00266015;
                12'd1502: logsin <= 24'd00266392;
                12'd1503: logsin <= 24'd00266769;
                12'd1504: logsin <= 24'd00267147;
                12'd1505: logsin <= 24'd00267525;
                12'd1506: logsin <= 24'd00267903;
                12'd1507: logsin <= 24'd00268281;
                12'd1508: logsin <= 24'd00268660;
                12'd1509: logsin <= 24'd00269039;
                12'd1510: logsin <= 24'd00269418;
                12'd1511: logsin <= 24'd00269798;
                12'd1512: logsin <= 24'd00270178;
                12'd1513: logsin <= 24'd00270558;
                12'd1514: logsin <= 24'd00270939;
                12'd1515: logsin <= 24'd00271319;
                12'd1516: logsin <= 24'd00271701;
                12'd1517: logsin <= 24'd00272082;
                12'd1518: logsin <= 24'd00272464;
                12'd1519: logsin <= 24'd00272846;
                12'd1520: logsin <= 24'd00273229;
                12'd1521: logsin <= 24'd00273612;
                12'd1522: logsin <= 24'd00273995;
                12'd1523: logsin <= 24'd00274378;
                12'd1524: logsin <= 24'd00274762;
                12'd1525: logsin <= 24'd00275146;
                12'd1526: logsin <= 24'd00275531;
                12'd1527: logsin <= 24'd00275915;
                12'd1528: logsin <= 24'd00276300;
                12'd1529: logsin <= 24'd00276686;
                12'd1530: logsin <= 24'd00277071;
                12'd1531: logsin <= 24'd00277458;
                12'd1532: logsin <= 24'd00277844;
                12'd1533: logsin <= 24'd00278231;
                12'd1534: logsin <= 24'd00278618;
                12'd1535: logsin <= 24'd00279005;
                12'd1536: logsin <= 24'd00279392;
                12'd1537: logsin <= 24'd00279780;
                12'd1538: logsin <= 24'd00280169;
                12'd1539: logsin <= 24'd00280557;
                12'd1540: logsin <= 24'd00280946;
                12'd1541: logsin <= 24'd00281336;
                12'd1542: logsin <= 24'd00281725;
                12'd1543: logsin <= 24'd00282115;
                12'd1544: logsin <= 24'd00282505;
                12'd1545: logsin <= 24'd00282896;
                12'd1546: logsin <= 24'd00283287;
                12'd1547: logsin <= 24'd00283678;
                12'd1548: logsin <= 24'd00284069;
                12'd1549: logsin <= 24'd00284461;
                12'd1550: logsin <= 24'd00284853;
                12'd1551: logsin <= 24'd00285246;
                12'd1552: logsin <= 24'd00285639;
                12'd1553: logsin <= 24'd00286032;
                12'd1554: logsin <= 24'd00286425;
                12'd1555: logsin <= 24'd00286819;
                12'd1556: logsin <= 24'd00287213;
                12'd1557: logsin <= 24'd00287608;
                12'd1558: logsin <= 24'd00288002;
                12'd1559: logsin <= 24'd00288397;
                12'd1560: logsin <= 24'd00288793;
                12'd1561: logsin <= 24'd00289188;
                12'd1562: logsin <= 24'd00289585;
                12'd1563: logsin <= 24'd00289981;
                12'd1564: logsin <= 24'd00290378;
                12'd1565: logsin <= 24'd00290775;
                12'd1566: logsin <= 24'd00291172;
                12'd1567: logsin <= 24'd00291570;
                12'd1568: logsin <= 24'd00291968;
                12'd1569: logsin <= 24'd00292366;
                12'd1570: logsin <= 24'd00292765;
                12'd1571: logsin <= 24'd00293164;
                12'd1572: logsin <= 24'd00293563;
                12'd1573: logsin <= 24'd00293963;
                12'd1574: logsin <= 24'd00294363;
                12'd1575: logsin <= 24'd00294763;
                12'd1576: logsin <= 24'd00295164;
                12'd1577: logsin <= 24'd00295565;
                12'd1578: logsin <= 24'd00295966;
                12'd1579: logsin <= 24'd00296368;
                12'd1580: logsin <= 24'd00296770;
                12'd1581: logsin <= 24'd00297172;
                12'd1582: logsin <= 24'd00297575;
                12'd1583: logsin <= 24'd00297977;
                12'd1584: logsin <= 24'd00298381;
                12'd1585: logsin <= 24'd00298784;
                12'd1586: logsin <= 24'd00299188;
                12'd1587: logsin <= 24'd00299593;
                12'd1588: logsin <= 24'd00299997;
                12'd1589: logsin <= 24'd00300402;
                12'd1590: logsin <= 24'd00300807;
                12'd1591: logsin <= 24'd00301213;
                12'd1592: logsin <= 24'd00301619;
                12'd1593: logsin <= 24'd00302025;
                12'd1594: logsin <= 24'd00302432;
                12'd1595: logsin <= 24'd00302839;
                12'd1596: logsin <= 24'd00303246;
                12'd1597: logsin <= 24'd00303654;
                12'd1598: logsin <= 24'd00304061;
                12'd1599: logsin <= 24'd00304470;
                12'd1600: logsin <= 24'd00304878;
                12'd1601: logsin <= 24'd00305287;
                12'd1602: logsin <= 24'd00305696;
                12'd1603: logsin <= 24'd00306106;
                12'd1604: logsin <= 24'd00306516;
                12'd1605: logsin <= 24'd00306926;
                12'd1606: logsin <= 24'd00307337;
                12'd1607: logsin <= 24'd00307748;
                12'd1608: logsin <= 24'd00308159;
                12'd1609: logsin <= 24'd00308571;
                12'd1610: logsin <= 24'd00308982;
                12'd1611: logsin <= 24'd00309395;
                12'd1612: logsin <= 24'd00309807;
                12'd1613: logsin <= 24'd00310220;
                12'd1614: logsin <= 24'd00310633;
                12'd1615: logsin <= 24'd00311047;
                12'd1616: logsin <= 24'd00311461;
                12'd1617: logsin <= 24'd00311875;
                12'd1618: logsin <= 24'd00312290;
                12'd1619: logsin <= 24'd00312705;
                12'd1620: logsin <= 24'd00313120;
                12'd1621: logsin <= 24'd00313536;
                12'd1622: logsin <= 24'd00313952;
                12'd1623: logsin <= 24'd00314368;
                12'd1624: logsin <= 24'd00314785;
                12'd1625: logsin <= 24'd00315201;
                12'd1626: logsin <= 24'd00315619;
                12'd1627: logsin <= 24'd00316036;
                12'd1628: logsin <= 24'd00316454;
                12'd1629: logsin <= 24'd00316873;
                12'd1630: logsin <= 24'd00317291;
                12'd1631: logsin <= 24'd00317710;
                12'd1632: logsin <= 24'd00318130;
                12'd1633: logsin <= 24'd00318549;
                12'd1634: logsin <= 24'd00318969;
                12'd1635: logsin <= 24'd00319390;
                12'd1636: logsin <= 24'd00319810;
                12'd1637: logsin <= 24'd00320231;
                12'd1638: logsin <= 24'd00320653;
                12'd1639: logsin <= 24'd00321074;
                12'd1640: logsin <= 24'd00321496;
                12'd1641: logsin <= 24'd00321919;
                12'd1642: logsin <= 24'd00322342;
                12'd1643: logsin <= 24'd00322765;
                12'd1644: logsin <= 24'd00323188;
                12'd1645: logsin <= 24'd00323612;
                12'd1646: logsin <= 24'd00324036;
                12'd1647: logsin <= 24'd00324460;
                12'd1648: logsin <= 24'd00324885;
                12'd1649: logsin <= 24'd00325310;
                12'd1650: logsin <= 24'd00325736;
                12'd1651: logsin <= 24'd00326161;
                12'd1652: logsin <= 24'd00326588;
                12'd1653: logsin <= 24'd00327014;
                12'd1654: logsin <= 24'd00327441;
                12'd1655: logsin <= 24'd00327868;
                12'd1656: logsin <= 24'd00328296;
                12'd1657: logsin <= 24'd00328723;
                12'd1658: logsin <= 24'd00329152;
                12'd1659: logsin <= 24'd00329580;
                12'd1660: logsin <= 24'd00330009;
                12'd1661: logsin <= 24'd00330438;
                12'd1662: logsin <= 24'd00330868;
                12'd1663: logsin <= 24'd00331298;
                12'd1664: logsin <= 24'd00331728;
                12'd1665: logsin <= 24'd00332159;
                12'd1666: logsin <= 24'd00332590;
                12'd1667: logsin <= 24'd00333021;
                12'd1668: logsin <= 24'd00333453;
                12'd1669: logsin <= 24'd00333885;
                12'd1670: logsin <= 24'd00334317;
                12'd1671: logsin <= 24'd00334750;
                12'd1672: logsin <= 24'd00335183;
                12'd1673: logsin <= 24'd00335616;
                12'd1674: logsin <= 24'd00336050;
                12'd1675: logsin <= 24'd00336484;
                12'd1676: logsin <= 24'd00336918;
                12'd1677: logsin <= 24'd00337353;
                12'd1678: logsin <= 24'd00337788;
                12'd1679: logsin <= 24'd00338223;
                12'd1680: logsin <= 24'd00338659;
                12'd1681: logsin <= 24'd00339095;
                12'd1682: logsin <= 24'd00339532;
                12'd1683: logsin <= 24'd00339969;
                12'd1684: logsin <= 24'd00340406;
                12'd1685: logsin <= 24'd00340844;
                12'd1686: logsin <= 24'd00341281;
                12'd1687: logsin <= 24'd00341720;
                12'd1688: logsin <= 24'd00342158;
                12'd1689: logsin <= 24'd00342597;
                12'd1690: logsin <= 24'd00343037;
                12'd1691: logsin <= 24'd00343476;
                12'd1692: logsin <= 24'd00343916;
                12'd1693: logsin <= 24'd00344357;
                12'd1694: logsin <= 24'd00344797;
                12'd1695: logsin <= 24'd00345238;
                12'd1696: logsin <= 24'd00345680;
                12'd1697: logsin <= 24'd00346121;
                12'd1698: logsin <= 24'd00346564;
                12'd1699: logsin <= 24'd00347006;
                12'd1700: logsin <= 24'd00347449;
                12'd1701: logsin <= 24'd00347892;
                12'd1702: logsin <= 24'd00348335;
                12'd1703: logsin <= 24'd00348779;
                12'd1704: logsin <= 24'd00349224;
                12'd1705: logsin <= 24'd00349668;
                12'd1706: logsin <= 24'd00350113;
                12'd1707: logsin <= 24'd00350558;
                12'd1708: logsin <= 24'd00351004;
                12'd1709: logsin <= 24'd00351450;
                12'd1710: logsin <= 24'd00351896;
                12'd1711: logsin <= 24'd00352343;
                12'd1712: logsin <= 24'd00352790;
                12'd1713: logsin <= 24'd00353237;
                12'd1714: logsin <= 24'd00353685;
                12'd1715: logsin <= 24'd00354133;
                12'd1716: logsin <= 24'd00354582;
                12'd1717: logsin <= 24'd00355031;
                12'd1718: logsin <= 24'd00355480;
                12'd1719: logsin <= 24'd00355929;
                12'd1720: logsin <= 24'd00356379;
                12'd1721: logsin <= 24'd00356829;
                12'd1722: logsin <= 24'd00357280;
                12'd1723: logsin <= 24'd00357731;
                12'd1724: logsin <= 24'd00358182;
                12'd1725: logsin <= 24'd00358634;
                12'd1726: logsin <= 24'd00359086;
                12'd1727: logsin <= 24'd00359538;
                12'd1728: logsin <= 24'd00359991;
                12'd1729: logsin <= 24'd00360444;
                12'd1730: logsin <= 24'd00360898;
                12'd1731: logsin <= 24'd00361352;
                12'd1732: logsin <= 24'd00361806;
                12'd1733: logsin <= 24'd00362260;
                12'd1734: logsin <= 24'd00362715;
                12'd1735: logsin <= 24'd00363170;
                12'd1736: logsin <= 24'd00363626;
                12'd1737: logsin <= 24'd00364082;
                12'd1738: logsin <= 24'd00364538;
                12'd1739: logsin <= 24'd00364995;
                12'd1740: logsin <= 24'd00365452;
                12'd1741: logsin <= 24'd00365909;
                12'd1742: logsin <= 24'd00366367;
                12'd1743: logsin <= 24'd00366825;
                12'd1744: logsin <= 24'd00367284;
                12'd1745: logsin <= 24'd00367743;
                12'd1746: logsin <= 24'd00368202;
                12'd1747: logsin <= 24'd00368662;
                12'd1748: logsin <= 24'd00369122;
                12'd1749: logsin <= 24'd00369582;
                12'd1750: logsin <= 24'd00370043;
                12'd1751: logsin <= 24'd00370504;
                12'd1752: logsin <= 24'd00370965;
                12'd1753: logsin <= 24'd00371427;
                12'd1754: logsin <= 24'd00371889;
                12'd1755: logsin <= 24'd00372351;
                12'd1756: logsin <= 24'd00372814;
                12'd1757: logsin <= 24'd00373277;
                12'd1758: logsin <= 24'd00373741;
                12'd1759: logsin <= 24'd00374205;
                12'd1760: logsin <= 24'd00374669;
                12'd1761: logsin <= 24'd00375134;
                12'd1762: logsin <= 24'd00375599;
                12'd1763: logsin <= 24'd00376064;
                12'd1764: logsin <= 24'd00376530;
                12'd1765: logsin <= 24'd00376996;
                12'd1766: logsin <= 24'd00377463;
                12'd1767: logsin <= 24'd00377930;
                12'd1768: logsin <= 24'd00378397;
                12'd1769: logsin <= 24'd00378865;
                12'd1770: logsin <= 24'd00379333;
                12'd1771: logsin <= 24'd00379801;
                12'd1772: logsin <= 24'd00380270;
                12'd1773: logsin <= 24'd00380739;
                12'd1774: logsin <= 24'd00381208;
                12'd1775: logsin <= 24'd00381678;
                12'd1776: logsin <= 24'd00382148;
                12'd1777: logsin <= 24'd00382619;
                12'd1778: logsin <= 24'd00383090;
                12'd1779: logsin <= 24'd00383561;
                12'd1780: logsin <= 24'd00384033;
                12'd1781: logsin <= 24'd00384505;
                12'd1782: logsin <= 24'd00384977;
                12'd1783: logsin <= 24'd00385450;
                12'd1784: logsin <= 24'd00385923;
                12'd1785: logsin <= 24'd00386396;
                12'd1786: logsin <= 24'd00386870;
                12'd1787: logsin <= 24'd00387345;
                12'd1788: logsin <= 24'd00387819;
                12'd1789: logsin <= 24'd00388294;
                12'd1790: logsin <= 24'd00388770;
                12'd1791: logsin <= 24'd00389245;
                12'd1792: logsin <= 24'd00389721;
                12'd1793: logsin <= 24'd00390198;
                12'd1794: logsin <= 24'd00390675;
                12'd1795: logsin <= 24'd00391152;
                12'd1796: logsin <= 24'd00391630;
                12'd1797: logsin <= 24'd00392107;
                12'd1798: logsin <= 24'd00392586;
                12'd1799: logsin <= 24'd00393065;
                12'd1800: logsin <= 24'd00393544;
                12'd1801: logsin <= 24'd00394023;
                12'd1802: logsin <= 24'd00394503;
                12'd1803: logsin <= 24'd00394983;
                12'd1804: logsin <= 24'd00395464;
                12'd1805: logsin <= 24'd00395945;
                12'd1806: logsin <= 24'd00396426;
                12'd1807: logsin <= 24'd00396908;
                12'd1808: logsin <= 24'd00397390;
                12'd1809: logsin <= 24'd00397872;
                12'd1810: logsin <= 24'd00398355;
                12'd1811: logsin <= 24'd00398838;
                12'd1812: logsin <= 24'd00399322;
                12'd1813: logsin <= 24'd00399806;
                12'd1814: logsin <= 24'd00400290;
                12'd1815: logsin <= 24'd00400775;
                12'd1816: logsin <= 24'd00401260;
                12'd1817: logsin <= 24'd00401746;
                12'd1818: logsin <= 24'd00402232;
                12'd1819: logsin <= 24'd00402718;
                12'd1820: logsin <= 24'd00403205;
                12'd1821: logsin <= 24'd00403692;
                12'd1822: logsin <= 24'd00404179;
                12'd1823: logsin <= 24'd00404667;
                12'd1824: logsin <= 24'd00405155;
                12'd1825: logsin <= 24'd00405643;
                12'd1826: logsin <= 24'd00406132;
                12'd1827: logsin <= 24'd00406622;
                12'd1828: logsin <= 24'd00407111;
                12'd1829: logsin <= 24'd00407601;
                12'd1830: logsin <= 24'd00408092;
                12'd1831: logsin <= 24'd00408583;
                12'd1832: logsin <= 24'd00409074;
                12'd1833: logsin <= 24'd00409565;
                12'd1834: logsin <= 24'd00410057;
                12'd1835: logsin <= 24'd00410550;
                12'd1836: logsin <= 24'd00411042;
                12'd1837: logsin <= 24'd00411535;
                12'd1838: logsin <= 24'd00412029;
                12'd1839: logsin <= 24'd00412523;
                12'd1840: logsin <= 24'd00413017;
                12'd1841: logsin <= 24'd00413512;
                12'd1842: logsin <= 24'd00414007;
                12'd1843: logsin <= 24'd00414502;
                12'd1844: logsin <= 24'd00414998;
                12'd1845: logsin <= 24'd00415494;
                12'd1846: logsin <= 24'd00415991;
                12'd1847: logsin <= 24'd00416488;
                12'd1848: logsin <= 24'd00416985;
                12'd1849: logsin <= 24'd00417483;
                12'd1850: logsin <= 24'd00417981;
                12'd1851: logsin <= 24'd00418479;
                12'd1852: logsin <= 24'd00418978;
                12'd1853: logsin <= 24'd00419477;
                12'd1854: logsin <= 24'd00419977;
                12'd1855: logsin <= 24'd00420477;
                12'd1856: logsin <= 24'd00420978;
                12'd1857: logsin <= 24'd00421478;
                12'd1858: logsin <= 24'd00421980;
                12'd1859: logsin <= 24'd00422481;
                12'd1860: logsin <= 24'd00422983;
                12'd1861: logsin <= 24'd00423486;
                12'd1862: logsin <= 24'd00423988;
                12'd1863: logsin <= 24'd00424491;
                12'd1864: logsin <= 24'd00424995;
                12'd1865: logsin <= 24'd00425499;
                12'd1866: logsin <= 24'd00426003;
                12'd1867: logsin <= 24'd00426508;
                12'd1868: logsin <= 24'd00427013;
                12'd1869: logsin <= 24'd00427519;
                12'd1870: logsin <= 24'd00428025;
                12'd1871: logsin <= 24'd00428531;
                12'd1872: logsin <= 24'd00429037;
                12'd1873: logsin <= 24'd00429545;
                12'd1874: logsin <= 24'd00430052;
                12'd1875: logsin <= 24'd00430560;
                12'd1876: logsin <= 24'd00431068;
                12'd1877: logsin <= 24'd00431577;
                12'd1878: logsin <= 24'd00432086;
                12'd1879: logsin <= 24'd00432595;
                12'd1880: logsin <= 24'd00433105;
                12'd1881: logsin <= 24'd00433615;
                12'd1882: logsin <= 24'd00434126;
                12'd1883: logsin <= 24'd00434637;
                12'd1884: logsin <= 24'd00435148;
                12'd1885: logsin <= 24'd00435660;
                12'd1886: logsin <= 24'd00436172;
                12'd1887: logsin <= 24'd00436685;
                12'd1888: logsin <= 24'd00437198;
                12'd1889: logsin <= 24'd00437711;
                12'd1890: logsin <= 24'd00438225;
                12'd1891: logsin <= 24'd00438739;
                12'd1892: logsin <= 24'd00439254;
                12'd1893: logsin <= 24'd00439769;
                12'd1894: logsin <= 24'd00440284;
                12'd1895: logsin <= 24'd00440800;
                12'd1896: logsin <= 24'd00441316;
                12'd1897: logsin <= 24'd00441833;
                12'd1898: logsin <= 24'd00442350;
                12'd1899: logsin <= 24'd00442867;
                12'd1900: logsin <= 24'd00443385;
                12'd1901: logsin <= 24'd00443903;
                12'd1902: logsin <= 24'd00444421;
                12'd1903: logsin <= 24'd00444940;
                12'd1904: logsin <= 24'd00445460;
                12'd1905: logsin <= 24'd00445979;
                12'd1906: logsin <= 24'd00446500;
                12'd1907: logsin <= 24'd00447020;
                12'd1908: logsin <= 24'd00447541;
                12'd1909: logsin <= 24'd00448063;
                12'd1910: logsin <= 24'd00448584;
                12'd1911: logsin <= 24'd00449106;
                12'd1912: logsin <= 24'd00449629;
                12'd1913: logsin <= 24'd00450152;
                12'd1914: logsin <= 24'd00450675;
                12'd1915: logsin <= 24'd00451199;
                12'd1916: logsin <= 24'd00451723;
                12'd1917: logsin <= 24'd00452248;
                12'd1918: logsin <= 24'd00452773;
                12'd1919: logsin <= 24'd00453298;
                12'd1920: logsin <= 24'd00453824;
                12'd1921: logsin <= 24'd00454350;
                12'd1922: logsin <= 24'd00454877;
                12'd1923: logsin <= 24'd00455404;
                12'd1924: logsin <= 24'd00455932;
                12'd1925: logsin <= 24'd00456459;
                12'd1926: logsin <= 24'd00456988;
                12'd1927: logsin <= 24'd00457516;
                12'd1928: logsin <= 24'd00458045;
                12'd1929: logsin <= 24'd00458575;
                12'd1930: logsin <= 24'd00459105;
                12'd1931: logsin <= 24'd00459635;
                12'd1932: logsin <= 24'd00460166;
                12'd1933: logsin <= 24'd00460697;
                12'd1934: logsin <= 24'd00461228;
                12'd1935: logsin <= 24'd00461760;
                12'd1936: logsin <= 24'd00462292;
                12'd1937: logsin <= 24'd00462825;
                12'd1938: logsin <= 24'd00463358;
                12'd1939: logsin <= 24'd00463892;
                12'd1940: logsin <= 24'd00464426;
                12'd1941: logsin <= 24'd00464960;
                12'd1942: logsin <= 24'd00465495;
                12'd1943: logsin <= 24'd00466030;
                12'd1944: logsin <= 24'd00466566;
                12'd1945: logsin <= 24'd00467102;
                12'd1946: logsin <= 24'd00467638;
                12'd1947: logsin <= 24'd00468175;
                12'd1948: logsin <= 24'd00468713;
                12'd1949: logsin <= 24'd00469250;
                12'd1950: logsin <= 24'd00469788;
                12'd1951: logsin <= 24'd00470327;
                12'd1952: logsin <= 24'd00470866;
                12'd1953: logsin <= 24'd00471405;
                12'd1954: logsin <= 24'd00471945;
                12'd1955: logsin <= 24'd00472485;
                12'd1956: logsin <= 24'd00473026;
                12'd1957: logsin <= 24'd00473567;
                12'd1958: logsin <= 24'd00474108;
                12'd1959: logsin <= 24'd00474650;
                12'd1960: logsin <= 24'd00475192;
                12'd1961: logsin <= 24'd00475735;
                12'd1962: logsin <= 24'd00476278;
                12'd1963: logsin <= 24'd00476821;
                12'd1964: logsin <= 24'd00477365;
                12'd1965: logsin <= 24'd00477910;
                12'd1966: logsin <= 24'd00478454;
                12'd1967: logsin <= 24'd00479000;
                12'd1968: logsin <= 24'd00479545;
                12'd1969: logsin <= 24'd00480091;
                12'd1970: logsin <= 24'd00480638;
                12'd1971: logsin <= 24'd00481184;
                12'd1972: logsin <= 24'd00481732;
                12'd1973: logsin <= 24'd00482279;
                12'd1974: logsin <= 24'd00482827;
                12'd1975: logsin <= 24'd00483376;
                12'd1976: logsin <= 24'd00483925;
                12'd1977: logsin <= 24'd00484474;
                12'd1978: logsin <= 24'd00485024;
                12'd1979: logsin <= 24'd00485574;
                12'd1980: logsin <= 24'd00486125;
                12'd1981: logsin <= 24'd00486676;
                12'd1982: logsin <= 24'd00487228;
                12'd1983: logsin <= 24'd00487780;
                12'd1984: logsin <= 24'd00488332;
                12'd1985: logsin <= 24'd00488885;
                12'd1986: logsin <= 24'd00489438;
                12'd1987: logsin <= 24'd00489991;
                12'd1988: logsin <= 24'd00490545;
                12'd1989: logsin <= 24'd00491100;
                12'd1990: logsin <= 24'd00491655;
                12'd1991: logsin <= 24'd00492210;
                12'd1992: logsin <= 24'd00492766;
                12'd1993: logsin <= 24'd00493322;
                12'd1994: logsin <= 24'd00493879;
                12'd1995: logsin <= 24'd00494436;
                12'd1996: logsin <= 24'd00494993;
                12'd1997: logsin <= 24'd00495551;
                12'd1998: logsin <= 24'd00496109;
                12'd1999: logsin <= 24'd00496668;
                12'd2000: logsin <= 24'd00497227;
                12'd2001: logsin <= 24'd00497787;
                12'd2002: logsin <= 24'd00498347;
                12'd2003: logsin <= 24'd00498907;
                12'd2004: logsin <= 24'd00499468;
                12'd2005: logsin <= 24'd00500030;
                12'd2006: logsin <= 24'd00500591;
                12'd2007: logsin <= 24'd00501153;
                12'd2008: logsin <= 24'd00501716;
                12'd2009: logsin <= 24'd00502279;
                12'd2010: logsin <= 24'd00502843;
                12'd2011: logsin <= 24'd00503406;
                12'd2012: logsin <= 24'd00503971;
                12'd2013: logsin <= 24'd00504536;
                12'd2014: logsin <= 24'd00505101;
                12'd2015: logsin <= 24'd00505666;
                12'd2016: logsin <= 24'd00506233;
                12'd2017: logsin <= 24'd00506799;
                12'd2018: logsin <= 24'd00507366;
                12'd2019: logsin <= 24'd00507933;
                12'd2020: logsin <= 24'd00508501;
                12'd2021: logsin <= 24'd00509069;
                12'd2022: logsin <= 24'd00509638;
                12'd2023: logsin <= 24'd00510207;
                12'd2024: logsin <= 24'd00510777;
                12'd2025: logsin <= 24'd00511347;
                12'd2026: logsin <= 24'd00511917;
                12'd2027: logsin <= 24'd00512488;
                12'd2028: logsin <= 24'd00513059;
                12'd2029: logsin <= 24'd00513631;
                12'd2030: logsin <= 24'd00514203;
                12'd2031: logsin <= 24'd00514776;
                12'd2032: logsin <= 24'd00515349;
                12'd2033: logsin <= 24'd00515923;
                12'd2034: logsin <= 24'd00516496;
                12'd2035: logsin <= 24'd00517071;
                12'd2036: logsin <= 24'd00517646;
                12'd2037: logsin <= 24'd00518221;
                12'd2038: logsin <= 24'd00518797;
                12'd2039: logsin <= 24'd00519373;
                12'd2040: logsin <= 24'd00519949;
                12'd2041: logsin <= 24'd00520526;
                12'd2042: logsin <= 24'd00521104;
                12'd2043: logsin <= 24'd00521682;
                12'd2044: logsin <= 24'd00522260;
                12'd2045: logsin <= 24'd00522839;
                12'd2046: logsin <= 24'd00523418;
                12'd2047: logsin <= 24'd00523998;
                12'd2048: logsin <= 24'd00524578;
                12'd2049: logsin <= 24'd00525159;
                12'd2050: logsin <= 24'd00525740;
                12'd2051: logsin <= 24'd00526321;
                12'd2052: logsin <= 24'd00526903;
                12'd2053: logsin <= 24'd00527486;
                12'd2054: logsin <= 24'd00528068;
                12'd2055: logsin <= 24'd00528652;
                12'd2056: logsin <= 24'd00529235;
                12'd2057: logsin <= 24'd00529819;
                12'd2058: logsin <= 24'd00530404;
                12'd2059: logsin <= 24'd00530989;
                12'd2060: logsin <= 24'd00531575;
                12'd2061: logsin <= 24'd00532161;
                12'd2062: logsin <= 24'd00532747;
                12'd2063: logsin <= 24'd00533334;
                12'd2064: logsin <= 24'd00533921;
                12'd2065: logsin <= 24'd00534509;
                12'd2066: logsin <= 24'd00535097;
                12'd2067: logsin <= 24'd00535686;
                12'd2068: logsin <= 24'd00536275;
                12'd2069: logsin <= 24'd00536864;
                12'd2070: logsin <= 24'd00537454;
                12'd2071: logsin <= 24'd00538045;
                12'd2072: logsin <= 24'd00538636;
                12'd2073: logsin <= 24'd00539227;
                12'd2074: logsin <= 24'd00539819;
                12'd2075: logsin <= 24'd00540411;
                12'd2076: logsin <= 24'd00541004;
                12'd2077: logsin <= 24'd00541597;
                12'd2078: logsin <= 24'd00542191;
                12'd2079: logsin <= 24'd00542785;
                12'd2080: logsin <= 24'd00543380;
                12'd2081: logsin <= 24'd00543975;
                12'd2082: logsin <= 24'd00544570;
                12'd2083: logsin <= 24'd00545166;
                12'd2084: logsin <= 24'd00545762;
                12'd2085: logsin <= 24'd00546359;
                12'd2086: logsin <= 24'd00546957;
                12'd2087: logsin <= 24'd00547554;
                12'd2088: logsin <= 24'd00548153;
                12'd2089: logsin <= 24'd00548751;
                12'd2090: logsin <= 24'd00549350;
                12'd2091: logsin <= 24'd00549950;
                12'd2092: logsin <= 24'd00550550;
                12'd2093: logsin <= 24'd00551151;
                12'd2094: logsin <= 24'd00551751;
                12'd2095: logsin <= 24'd00552353;
                12'd2096: logsin <= 24'd00552955;
                12'd2097: logsin <= 24'd00553557;
                12'd2098: logsin <= 24'd00554160;
                12'd2099: logsin <= 24'd00554763;
                12'd2100: logsin <= 24'd00555367;
                12'd2101: logsin <= 24'd00555971;
                12'd2102: logsin <= 24'd00556576;
                12'd2103: logsin <= 24'd00557181;
                12'd2104: logsin <= 24'd00557787;
                12'd2105: logsin <= 24'd00558393;
                12'd2106: logsin <= 24'd00558999;
                12'd2107: logsin <= 24'd00559606;
                12'd2108: logsin <= 24'd00560214;
                12'd2109: logsin <= 24'd00560822;
                12'd2110: logsin <= 24'd00561430;
                12'd2111: logsin <= 24'd00562039;
                12'd2112: logsin <= 24'd00562648;
                12'd2113: logsin <= 24'd00563258;
                12'd2114: logsin <= 24'd00563868;
                12'd2115: logsin <= 24'd00564479;
                12'd2116: logsin <= 24'd00565090;
                12'd2117: logsin <= 24'd00565702;
                12'd2118: logsin <= 24'd00566314;
                12'd2119: logsin <= 24'd00566927;
                12'd2120: logsin <= 24'd00567540;
                12'd2121: logsin <= 24'd00568154;
                12'd2122: logsin <= 24'd00568768;
                12'd2123: logsin <= 24'd00569382;
                12'd2124: logsin <= 24'd00569997;
                12'd2125: logsin <= 24'd00570613;
                12'd2126: logsin <= 24'd00571229;
                12'd2127: logsin <= 24'd00571845;
                12'd2128: logsin <= 24'd00572462;
                12'd2129: logsin <= 24'd00573079;
                12'd2130: logsin <= 24'd00573697;
                12'd2131: logsin <= 24'd00574315;
                12'd2132: logsin <= 24'd00574934;
                12'd2133: logsin <= 24'd00575553;
                12'd2134: logsin <= 24'd00576173;
                12'd2135: logsin <= 24'd00576793;
                12'd2136: logsin <= 24'd00577414;
                12'd2137: logsin <= 24'd00578035;
                12'd2138: logsin <= 24'd00578657;
                12'd2139: logsin <= 24'd00579279;
                12'd2140: logsin <= 24'd00579901;
                12'd2141: logsin <= 24'd00580525;
                12'd2142: logsin <= 24'd00581148;
                12'd2143: logsin <= 24'd00581772;
                12'd2144: logsin <= 24'd00582397;
                12'd2145: logsin <= 24'd00583022;
                12'd2146: logsin <= 24'd00583647;
                12'd2147: logsin <= 24'd00584273;
                12'd2148: logsin <= 24'd00584899;
                12'd2149: logsin <= 24'd00585526;
                12'd2150: logsin <= 24'd00586154;
                12'd2151: logsin <= 24'd00586782;
                12'd2152: logsin <= 24'd00587410;
                12'd2153: logsin <= 24'd00588039;
                12'd2154: logsin <= 24'd00588668;
                12'd2155: logsin <= 24'd00589298;
                12'd2156: logsin <= 24'd00589928;
                12'd2157: logsin <= 24'd00590559;
                12'd2158: logsin <= 24'd00591190;
                12'd2159: logsin <= 24'd00591822;
                12'd2160: logsin <= 24'd00592454;
                12'd2161: logsin <= 24'd00593087;
                12'd2162: logsin <= 24'd00593720;
                12'd2163: logsin <= 24'd00594354;
                12'd2164: logsin <= 24'd00594988;
                12'd2165: logsin <= 24'd00595623;
                12'd2166: logsin <= 24'd00596258;
                12'd2167: logsin <= 24'd00596894;
                12'd2168: logsin <= 24'd00597530;
                12'd2169: logsin <= 24'd00598167;
                12'd2170: logsin <= 24'd00598804;
                12'd2171: logsin <= 24'd00599441;
                12'd2172: logsin <= 24'd00600079;
                12'd2173: logsin <= 24'd00600718;
                12'd2174: logsin <= 24'd00601357;
                12'd2175: logsin <= 24'd00601997;
                12'd2176: logsin <= 24'd00602637;
                12'd2177: logsin <= 24'd00603277;
                12'd2178: logsin <= 24'd00603919;
                12'd2179: logsin <= 24'd00604560;
                12'd2180: logsin <= 24'd00605202;
                12'd2181: logsin <= 24'd00605845;
                12'd2182: logsin <= 24'd00606488;
                12'd2183: logsin <= 24'd00607131;
                12'd2184: logsin <= 24'd00607775;
                12'd2185: logsin <= 24'd00608420;
                12'd2186: logsin <= 24'd00609065;
                12'd2187: logsin <= 24'd00609711;
                12'd2188: logsin <= 24'd00610357;
                12'd2189: logsin <= 24'd00611003;
                12'd2190: logsin <= 24'd00611650;
                12'd2191: logsin <= 24'd00612298;
                12'd2192: logsin <= 24'd00612946;
                12'd2193: logsin <= 24'd00613594;
                12'd2194: logsin <= 24'd00614243;
                12'd2195: logsin <= 24'd00614893;
                12'd2196: logsin <= 24'd00615543;
                12'd2197: logsin <= 24'd00616193;
                12'd2198: logsin <= 24'd00616844;
                12'd2199: logsin <= 24'd00617496;
                12'd2200: logsin <= 24'd00618148;
                12'd2201: logsin <= 24'd00618801;
                12'd2202: logsin <= 24'd00619454;
                12'd2203: logsin <= 24'd00620107;
                12'd2204: logsin <= 24'd00620761;
                12'd2205: logsin <= 24'd00621416;
                12'd2206: logsin <= 24'd00622071;
                12'd2207: logsin <= 24'd00622727;
                12'd2208: logsin <= 24'd00623383;
                12'd2209: logsin <= 24'd00624039;
                12'd2210: logsin <= 24'd00624696;
                12'd2211: logsin <= 24'd00625354;
                12'd2212: logsin <= 24'd00626012;
                12'd2213: logsin <= 24'd00626671;
                12'd2214: logsin <= 24'd00627330;
                12'd2215: logsin <= 24'd00627989;
                12'd2216: logsin <= 24'd00628650;
                12'd2217: logsin <= 24'd00629310;
                12'd2218: logsin <= 24'd00629971;
                12'd2219: logsin <= 24'd00630633;
                12'd2220: logsin <= 24'd00631295;
                12'd2221: logsin <= 24'd00631958;
                12'd2222: logsin <= 24'd00632621;
                12'd2223: logsin <= 24'd00633285;
                12'd2224: logsin <= 24'd00633949;
                12'd2225: logsin <= 24'd00634614;
                12'd2226: logsin <= 24'd00635279;
                12'd2227: logsin <= 24'd00635945;
                12'd2228: logsin <= 24'd00636612;
                12'd2229: logsin <= 24'd00637278;
                12'd2230: logsin <= 24'd00637946;
                12'd2231: logsin <= 24'd00638614;
                12'd2232: logsin <= 24'd00639282;
                12'd2233: logsin <= 24'd00639951;
                12'd2234: logsin <= 24'd00640620;
                12'd2235: logsin <= 24'd00641290;
                12'd2236: logsin <= 24'd00641961;
                12'd2237: logsin <= 24'd00642632;
                12'd2238: logsin <= 24'd00643303;
                12'd2239: logsin <= 24'd00643975;
                12'd2240: logsin <= 24'd00644648;
                12'd2241: logsin <= 24'd00645321;
                12'd2242: logsin <= 24'd00645994;
                12'd2243: logsin <= 24'd00646669;
                12'd2244: logsin <= 24'd00647343;
                12'd2245: logsin <= 24'd00648018;
                12'd2246: logsin <= 24'd00648694;
                12'd2247: logsin <= 24'd00649370;
                12'd2248: logsin <= 24'd00650047;
                12'd2249: logsin <= 24'd00650724;
                12'd2250: logsin <= 24'd00651402;
                12'd2251: logsin <= 24'd00652080;
                12'd2252: logsin <= 24'd00652759;
                12'd2253: logsin <= 24'd00653439;
                12'd2254: logsin <= 24'd00654118;
                12'd2255: logsin <= 24'd00654799;
                12'd2256: logsin <= 24'd00655480;
                12'd2257: logsin <= 24'd00656161;
                12'd2258: logsin <= 24'd00656843;
                12'd2259: logsin <= 24'd00657526;
                12'd2260: logsin <= 24'd00658209;
                12'd2261: logsin <= 24'd00658892;
                12'd2262: logsin <= 24'd00659577;
                12'd2263: logsin <= 24'd00660261;
                12'd2264: logsin <= 24'd00660946;
                12'd2265: logsin <= 24'd00661632;
                12'd2266: logsin <= 24'd00662318;
                12'd2267: logsin <= 24'd00663005;
                12'd2268: logsin <= 24'd00663693;
                12'd2269: logsin <= 24'd00664380;
                12'd2270: logsin <= 24'd00665069;
                12'd2271: logsin <= 24'd00665758;
                12'd2272: logsin <= 24'd00666447;
                12'd2273: logsin <= 24'd00667137;
                12'd2274: logsin <= 24'd00667828;
                12'd2275: logsin <= 24'd00668519;
                12'd2276: logsin <= 24'd00669211;
                12'd2277: logsin <= 24'd00669903;
                12'd2278: logsin <= 24'd00670595;
                12'd2279: logsin <= 24'd00671289;
                12'd2280: logsin <= 24'd00671982;
                12'd2281: logsin <= 24'd00672677;
                12'd2282: logsin <= 24'd00673372;
                12'd2283: logsin <= 24'd00674067;
                12'd2284: logsin <= 24'd00674763;
                12'd2285: logsin <= 24'd00675460;
                12'd2286: logsin <= 24'd00676157;
                12'd2287: logsin <= 24'd00676854;
                12'd2288: logsin <= 24'd00677552;
                12'd2289: logsin <= 24'd00678251;
                12'd2290: logsin <= 24'd00678950;
                12'd2291: logsin <= 24'd00679650;
                12'd2292: logsin <= 24'd00680350;
                12'd2293: logsin <= 24'd00681051;
                12'd2294: logsin <= 24'd00681752;
                12'd2295: logsin <= 24'd00682454;
                12'd2296: logsin <= 24'd00683157;
                12'd2297: logsin <= 24'd00683860;
                12'd2298: logsin <= 24'd00684564;
                12'd2299: logsin <= 24'd00685268;
                12'd2300: logsin <= 24'd00685972;
                12'd2301: logsin <= 24'd00686678;
                12'd2302: logsin <= 24'd00687383;
                12'd2303: logsin <= 24'd00688090;
                12'd2304: logsin <= 24'd00688797;
                12'd2305: logsin <= 24'd00689504;
                12'd2306: logsin <= 24'd00690212;
                12'd2307: logsin <= 24'd00690921;
                12'd2308: logsin <= 24'd00691630;
                12'd2309: logsin <= 24'd00692340;
                12'd2310: logsin <= 24'd00693050;
                12'd2311: logsin <= 24'd00693761;
                12'd2312: logsin <= 24'd00694472;
                12'd2313: logsin <= 24'd00695184;
                12'd2314: logsin <= 24'd00695896;
                12'd2315: logsin <= 24'd00696609;
                12'd2316: logsin <= 24'd00697323;
                12'd2317: logsin <= 24'd00698037;
                12'd2318: logsin <= 24'd00698752;
                12'd2319: logsin <= 24'd00699467;
                12'd2320: logsin <= 24'd00700183;
                12'd2321: logsin <= 24'd00700899;
                12'd2322: logsin <= 24'd00701616;
                12'd2323: logsin <= 24'd00702334;
                12'd2324: logsin <= 24'd00703052;
                12'd2325: logsin <= 24'd00703770;
                12'd2326: logsin <= 24'd00704489;
                12'd2327: logsin <= 24'd00705209;
                12'd2328: logsin <= 24'd00705930;
                12'd2329: logsin <= 24'd00706650;
                12'd2330: logsin <= 24'd00707372;
                12'd2331: logsin <= 24'd00708094;
                12'd2332: logsin <= 24'd00708817;
                12'd2333: logsin <= 24'd00709540;
                12'd2334: logsin <= 24'd00710263;
                12'd2335: logsin <= 24'd00710988;
                12'd2336: logsin <= 24'd00711713;
                12'd2337: logsin <= 24'd00712438;
                12'd2338: logsin <= 24'd00713164;
                12'd2339: logsin <= 24'd00713891;
                12'd2340: logsin <= 24'd00714618;
                12'd2341: logsin <= 24'd00715345;
                12'd2342: logsin <= 24'd00716074;
                12'd2343: logsin <= 24'd00716803;
                12'd2344: logsin <= 24'd00717532;
                12'd2345: logsin <= 24'd00718262;
                12'd2346: logsin <= 24'd00718993;
                12'd2347: logsin <= 24'd00719724;
                12'd2348: logsin <= 24'd00720456;
                12'd2349: logsin <= 24'd00721188;
                12'd2350: logsin <= 24'd00721921;
                12'd2351: logsin <= 24'd00722654;
                12'd2352: logsin <= 24'd00723388;
                12'd2353: logsin <= 24'd00724123;
                12'd2354: logsin <= 24'd00724858;
                12'd2355: logsin <= 24'd00725594;
                12'd2356: logsin <= 24'd00726330;
                12'd2357: logsin <= 24'd00727067;
                12'd2358: logsin <= 24'd00727805;
                12'd2359: logsin <= 24'd00728543;
                12'd2360: logsin <= 24'd00729282;
                12'd2361: logsin <= 24'd00730021;
                12'd2362: logsin <= 24'd00730761;
                12'd2363: logsin <= 24'd00731501;
                12'd2364: logsin <= 24'd00732242;
                12'd2365: logsin <= 24'd00732984;
                12'd2366: logsin <= 24'd00733726;
                12'd2367: logsin <= 24'd00734469;
                12'd2368: logsin <= 24'd00735212;
                12'd2369: logsin <= 24'd00735956;
                12'd2370: logsin <= 24'd00736701;
                12'd2371: logsin <= 24'd00737446;
                12'd2372: logsin <= 24'd00738192;
                12'd2373: logsin <= 24'd00738938;
                12'd2374: logsin <= 24'd00739685;
                12'd2375: logsin <= 24'd00740432;
                12'd2376: logsin <= 24'd00741181;
                12'd2377: logsin <= 24'd00741929;
                12'd2378: logsin <= 24'd00742679;
                12'd2379: logsin <= 24'd00743428;
                12'd2380: logsin <= 24'd00744179;
                12'd2381: logsin <= 24'd00744930;
                12'd2382: logsin <= 24'd00745682;
                12'd2383: logsin <= 24'd00746434;
                12'd2384: logsin <= 24'd00747187;
                12'd2385: logsin <= 24'd00747940;
                12'd2386: logsin <= 24'd00748694;
                12'd2387: logsin <= 24'd00749449;
                12'd2388: logsin <= 24'd00750204;
                12'd2389: logsin <= 24'd00750960;
                12'd2390: logsin <= 24'd00751717;
                12'd2391: logsin <= 24'd00752474;
                12'd2392: logsin <= 24'd00753231;
                12'd2393: logsin <= 24'd00753989;
                12'd2394: logsin <= 24'd00754748;
                12'd2395: logsin <= 24'd00755508;
                12'd2396: logsin <= 24'd00756268;
                12'd2397: logsin <= 24'd00757029;
                12'd2398: logsin <= 24'd00757790;
                12'd2399: logsin <= 24'd00758552;
                12'd2400: logsin <= 24'd00759314;
                12'd2401: logsin <= 24'd00760077;
                12'd2402: logsin <= 24'd00760841;
                12'd2403: logsin <= 24'd00761605;
                12'd2404: logsin <= 24'd00762370;
                12'd2405: logsin <= 24'd00763136;
                12'd2406: logsin <= 24'd00763902;
                12'd2407: logsin <= 24'd00764669;
                12'd2408: logsin <= 24'd00765436;
                12'd2409: logsin <= 24'd00766204;
                12'd2410: logsin <= 24'd00766973;
                12'd2411: logsin <= 24'd00767742;
                12'd2412: logsin <= 24'd00768512;
                12'd2413: logsin <= 24'd00769282;
                12'd2414: logsin <= 24'd00770053;
                12'd2415: logsin <= 24'd00770825;
                12'd2416: logsin <= 24'd00771597;
                12'd2417: logsin <= 24'd00772370;
                12'd2418: logsin <= 24'd00773144;
                12'd2419: logsin <= 24'd00773918;
                12'd2420: logsin <= 24'd00774692;
                12'd2421: logsin <= 24'd00775468;
                12'd2422: logsin <= 24'd00776244;
                12'd2423: logsin <= 24'd00777020;
                12'd2424: logsin <= 24'd00777798;
                12'd2425: logsin <= 24'd00778576;
                12'd2426: logsin <= 24'd00779354;
                12'd2427: logsin <= 24'd00780133;
                12'd2428: logsin <= 24'd00780913;
                12'd2429: logsin <= 24'd00781693;
                12'd2430: logsin <= 24'd00782474;
                12'd2431: logsin <= 24'd00783256;
                12'd2432: logsin <= 24'd00784038;
                12'd2433: logsin <= 24'd00784821;
                12'd2434: logsin <= 24'd00785604;
                12'd2435: logsin <= 24'd00786388;
                12'd2436: logsin <= 24'd00787173;
                12'd2437: logsin <= 24'd00787959;
                12'd2438: logsin <= 24'd00788745;
                12'd2439: logsin <= 24'd00789531;
                12'd2440: logsin <= 24'd00790318;
                12'd2441: logsin <= 24'd00791106;
                12'd2442: logsin <= 24'd00791895;
                12'd2443: logsin <= 24'd00792684;
                12'd2444: logsin <= 24'd00793474;
                12'd2445: logsin <= 24'd00794264;
                12'd2446: logsin <= 24'd00795055;
                12'd2447: logsin <= 24'd00795847;
                12'd2448: logsin <= 24'd00796639;
                12'd2449: logsin <= 24'd00797432;
                12'd2450: logsin <= 24'd00798226;
                12'd2451: logsin <= 24'd00799020;
                12'd2452: logsin <= 24'd00799815;
                12'd2453: logsin <= 24'd00800611;
                12'd2454: logsin <= 24'd00801407;
                12'd2455: logsin <= 24'd00802204;
                12'd2456: logsin <= 24'd00803001;
                12'd2457: logsin <= 24'd00803799;
                12'd2458: logsin <= 24'd00804598;
                12'd2459: logsin <= 24'd00805397;
                12'd2460: logsin <= 24'd00806198;
                12'd2461: logsin <= 24'd00806998;
                12'd2462: logsin <= 24'd00807800;
                12'd2463: logsin <= 24'd00808602;
                12'd2464: logsin <= 24'd00809404;
                12'd2465: logsin <= 24'd00810207;
                12'd2466: logsin <= 24'd00811011;
                12'd2467: logsin <= 24'd00811816;
                12'd2468: logsin <= 24'd00812621;
                12'd2469: logsin <= 24'd00813427;
                12'd2470: logsin <= 24'd00814234;
                12'd2471: logsin <= 24'd00815041;
                12'd2472: logsin <= 24'd00815849;
                12'd2473: logsin <= 24'd00816657;
                12'd2474: logsin <= 24'd00817466;
                12'd2475: logsin <= 24'd00818276;
                12'd2476: logsin <= 24'd00819087;
                12'd2477: logsin <= 24'd00819898;
                12'd2478: logsin <= 24'd00820709;
                12'd2479: logsin <= 24'd00821522;
                12'd2480: logsin <= 24'd00822335;
                12'd2481: logsin <= 24'd00823149;
                12'd2482: logsin <= 24'd00823963;
                12'd2483: logsin <= 24'd00824778;
                12'd2484: logsin <= 24'd00825594;
                12'd2485: logsin <= 24'd00826410;
                12'd2486: logsin <= 24'd00827227;
                12'd2487: logsin <= 24'd00828045;
                12'd2488: logsin <= 24'd00828864;
                12'd2489: logsin <= 24'd00829683;
                12'd2490: logsin <= 24'd00830502;
                12'd2491: logsin <= 24'd00831323;
                12'd2492: logsin <= 24'd00832144;
                12'd2493: logsin <= 24'd00832966;
                12'd2494: logsin <= 24'd00833788;
                12'd2495: logsin <= 24'd00834611;
                12'd2496: logsin <= 24'd00835435;
                12'd2497: logsin <= 24'd00836259;
                12'd2498: logsin <= 24'd00837084;
                12'd2499: logsin <= 24'd00837910;
                12'd2500: logsin <= 24'd00838736;
                12'd2501: logsin <= 24'd00839564;
                12'd2502: logsin <= 24'd00840391;
                12'd2503: logsin <= 24'd00841220;
                12'd2504: logsin <= 24'd00842049;
                12'd2505: logsin <= 24'd00842879;
                12'd2506: logsin <= 24'd00843709;
                12'd2507: logsin <= 24'd00844540;
                12'd2508: logsin <= 24'd00845372;
                12'd2509: logsin <= 24'd00846205;
                12'd2510: logsin <= 24'd00847038;
                12'd2511: logsin <= 24'd00847872;
                12'd2512: logsin <= 24'd00848706;
                12'd2513: logsin <= 24'd00849542;
                12'd2514: logsin <= 24'd00850378;
                12'd2515: logsin <= 24'd00851214;
                12'd2516: logsin <= 24'd00852051;
                12'd2517: logsin <= 24'd00852889;
                12'd2518: logsin <= 24'd00853728;
                12'd2519: logsin <= 24'd00854568;
                12'd2520: logsin <= 24'd00855408;
                12'd2521: logsin <= 24'd00856248;
                12'd2522: logsin <= 24'd00857090;
                12'd2523: logsin <= 24'd00857932;
                12'd2524: logsin <= 24'd00858775;
                12'd2525: logsin <= 24'd00859618;
                12'd2526: logsin <= 24'd00860462;
                12'd2527: logsin <= 24'd00861307;
                12'd2528: logsin <= 24'd00862153;
                12'd2529: logsin <= 24'd00862999;
                12'd2530: logsin <= 24'd00863846;
                12'd2531: logsin <= 24'd00864694;
                12'd2532: logsin <= 24'd00865542;
                12'd2533: logsin <= 24'd00866391;
                12'd2534: logsin <= 24'd00867241;
                12'd2535: logsin <= 24'd00868092;
                12'd2536: logsin <= 24'd00868943;
                12'd2537: logsin <= 24'd00869795;
                12'd2538: logsin <= 24'd00870647;
                12'd2539: logsin <= 24'd00871501;
                12'd2540: logsin <= 24'd00872355;
                12'd2541: logsin <= 24'd00873209;
                12'd2542: logsin <= 24'd00874065;
                12'd2543: logsin <= 24'd00874921;
                12'd2544: logsin <= 24'd00875778;
                12'd2545: logsin <= 24'd00876635;
                12'd2546: logsin <= 24'd00877493;
                12'd2547: logsin <= 24'd00878352;
                12'd2548: logsin <= 24'd00879212;
                12'd2549: logsin <= 24'd00880072;
                12'd2550: logsin <= 24'd00880933;
                12'd2551: logsin <= 24'd00881795;
                12'd2552: logsin <= 24'd00882658;
                12'd2553: logsin <= 24'd00883521;
                12'd2554: logsin <= 24'd00884385;
                12'd2555: logsin <= 24'd00885249;
                12'd2556: logsin <= 24'd00886115;
                12'd2557: logsin <= 24'd00886981;
                12'd2558: logsin <= 24'd00887848;
                12'd2559: logsin <= 24'd00888715;
                12'd2560: logsin <= 24'd00889583;
                12'd2561: logsin <= 24'd00890452;
                12'd2562: logsin <= 24'd00891322;
                12'd2563: logsin <= 24'd00892193;
                12'd2564: logsin <= 24'd00893064;
                12'd2565: logsin <= 24'd00893936;
                12'd2566: logsin <= 24'd00894808;
                12'd2567: logsin <= 24'd00895681;
                12'd2568: logsin <= 24'd00896555;
                12'd2569: logsin <= 24'd00897430;
                12'd2570: logsin <= 24'd00898306;
                12'd2571: logsin <= 24'd00899182;
                12'd2572: logsin <= 24'd00900059;
                12'd2573: logsin <= 24'd00900937;
                12'd2574: logsin <= 24'd00901815;
                12'd2575: logsin <= 24'd00902694;
                12'd2576: logsin <= 24'd00903574;
                12'd2577: logsin <= 24'd00904455;
                12'd2578: logsin <= 24'd00905336;
                12'd2579: logsin <= 24'd00906218;
                12'd2580: logsin <= 24'd00907101;
                12'd2581: logsin <= 24'd00907984;
                12'd2582: logsin <= 24'd00908869;
                12'd2583: logsin <= 24'd00909754;
                12'd2584: logsin <= 24'd00910640;
                12'd2585: logsin <= 24'd00911526;
                12'd2586: logsin <= 24'd00912413;
                12'd2587: logsin <= 24'd00913301;
                12'd2588: logsin <= 24'd00914190;
                12'd2589: logsin <= 24'd00915080;
                12'd2590: logsin <= 24'd00915970;
                12'd2591: logsin <= 24'd00916861;
                12'd2592: logsin <= 24'd00917753;
                12'd2593: logsin <= 24'd00918645;
                12'd2594: logsin <= 24'd00919538;
                12'd2595: logsin <= 24'd00920432;
                12'd2596: logsin <= 24'd00921327;
                12'd2597: logsin <= 24'd00922223;
                12'd2598: logsin <= 24'd00923119;
                12'd2599: logsin <= 24'd00924016;
                12'd2600: logsin <= 24'd00924914;
                12'd2601: logsin <= 24'd00925812;
                12'd2602: logsin <= 24'd00926711;
                12'd2603: logsin <= 24'd00927611;
                12'd2604: logsin <= 24'd00928512;
                12'd2605: logsin <= 24'd00929414;
                12'd2606: logsin <= 24'd00930316;
                12'd2607: logsin <= 24'd00931219;
                12'd2608: logsin <= 24'd00932123;
                12'd2609: logsin <= 24'd00933028;
                12'd2610: logsin <= 24'd00933933;
                12'd2611: logsin <= 24'd00934839;
                12'd2612: logsin <= 24'd00935746;
                12'd2613: logsin <= 24'd00936654;
                12'd2614: logsin <= 24'd00937562;
                12'd2615: logsin <= 24'd00938471;
                12'd2616: logsin <= 24'd00939381;
                12'd2617: logsin <= 24'd00940292;
                12'd2618: logsin <= 24'd00941203;
                12'd2619: logsin <= 24'd00942116;
                12'd2620: logsin <= 24'd00943029;
                12'd2621: logsin <= 24'd00943942;
                12'd2622: logsin <= 24'd00944857;
                12'd2623: logsin <= 24'd00945772;
                12'd2624: logsin <= 24'd00946689;
                12'd2625: logsin <= 24'd00947605;
                12'd2626: logsin <= 24'd00948523;
                12'd2627: logsin <= 24'd00949442;
                12'd2628: logsin <= 24'd00950361;
                12'd2629: logsin <= 24'd00951281;
                12'd2630: logsin <= 24'd00952202;
                12'd2631: logsin <= 24'd00953123;
                12'd2632: logsin <= 24'd00954046;
                12'd2633: logsin <= 24'd00954969;
                12'd2634: logsin <= 24'd00955893;
                12'd2635: logsin <= 24'd00956818;
                12'd2636: logsin <= 24'd00957743;
                12'd2637: logsin <= 24'd00958670;
                12'd2638: logsin <= 24'd00959597;
                12'd2639: logsin <= 24'd00960525;
                12'd2640: logsin <= 24'd00961453;
                12'd2641: logsin <= 24'd00962383;
                12'd2642: logsin <= 24'd00963313;
                12'd2643: logsin <= 24'd00964244;
                12'd2644: logsin <= 24'd00965176;
                12'd2645: logsin <= 24'd00966109;
                12'd2646: logsin <= 24'd00967042;
                12'd2647: logsin <= 24'd00967976;
                12'd2648: logsin <= 24'd00968912;
                12'd2649: logsin <= 24'd00969847;
                12'd2650: logsin <= 24'd00970784;
                12'd2651: logsin <= 24'd00971722;
                12'd2652: logsin <= 24'd00972660;
                12'd2653: logsin <= 24'd00973599;
                12'd2654: logsin <= 24'd00974539;
                12'd2655: logsin <= 24'd00975480;
                12'd2656: logsin <= 24'd00976421;
                12'd2657: logsin <= 24'd00977363;
                12'd2658: logsin <= 24'd00978307;
                12'd2659: logsin <= 24'd00979250;
                12'd2660: logsin <= 24'd00980195;
                12'd2661: logsin <= 24'd00981141;
                12'd2662: logsin <= 24'd00982087;
                12'd2663: logsin <= 24'd00983034;
                12'd2664: logsin <= 24'd00983982;
                12'd2665: logsin <= 24'd00984931;
                12'd2666: logsin <= 24'd00985881;
                12'd2667: logsin <= 24'd00986831;
                12'd2668: logsin <= 24'd00987783;
                12'd2669: logsin <= 24'd00988735;
                12'd2670: logsin <= 24'd00989688;
                12'd2671: logsin <= 24'd00990641;
                12'd2672: logsin <= 24'd00991596;
                12'd2673: logsin <= 24'd00992551;
                12'd2674: logsin <= 24'd00993508;
                12'd2675: logsin <= 24'd00994465;
                12'd2676: logsin <= 24'd00995423;
                12'd2677: logsin <= 24'd00996381;
                12'd2678: logsin <= 24'd00997341;
                12'd2679: logsin <= 24'd00998301;
                12'd2680: logsin <= 24'd00999262;
                12'd2681: logsin <= 24'd01000224;
                12'd2682: logsin <= 24'd01001187;
                12'd2683: logsin <= 24'd01002151;
                12'd2684: logsin <= 24'd01003116;
                12'd2685: logsin <= 24'd01004081;
                12'd2686: logsin <= 24'd01005047;
                12'd2687: logsin <= 24'd01006014;
                12'd2688: logsin <= 24'd01006982;
                12'd2689: logsin <= 24'd01007951;
                12'd2690: logsin <= 24'd01008920;
                12'd2691: logsin <= 24'd01009891;
                12'd2692: logsin <= 24'd01010862;
                12'd2693: logsin <= 24'd01011834;
                12'd2694: logsin <= 24'd01012807;
                12'd2695: logsin <= 24'd01013781;
                12'd2696: logsin <= 24'd01014756;
                12'd2697: logsin <= 24'd01015731;
                12'd2698: logsin <= 24'd01016708;
                12'd2699: logsin <= 24'd01017685;
                12'd2700: logsin <= 24'd01018663;
                12'd2701: logsin <= 24'd01019642;
                12'd2702: logsin <= 24'd01020622;
                12'd2703: logsin <= 24'd01021602;
                12'd2704: logsin <= 24'd01022584;
                12'd2705: logsin <= 24'd01023566;
                12'd2706: logsin <= 24'd01024550;
                12'd2707: logsin <= 24'd01025534;
                12'd2708: logsin <= 24'd01026519;
                12'd2709: logsin <= 24'd01027504;
                12'd2710: logsin <= 24'd01028491;
                12'd2711: logsin <= 24'd01029479;
                12'd2712: logsin <= 24'd01030467;
                12'd2713: logsin <= 24'd01031456;
                12'd2714: logsin <= 24'd01032447;
                12'd2715: logsin <= 24'd01033438;
                12'd2716: logsin <= 24'd01034430;
                12'd2717: logsin <= 24'd01035422;
                12'd2718: logsin <= 24'd01036416;
                12'd2719: logsin <= 24'd01037411;
                12'd2720: logsin <= 24'd01038406;
                12'd2721: logsin <= 24'd01039402;
                12'd2722: logsin <= 24'd01040399;
                12'd2723: logsin <= 24'd01041397;
                12'd2724: logsin <= 24'd01042396;
                12'd2725: logsin <= 24'd01043396;
                12'd2726: logsin <= 24'd01044397;
                12'd2727: logsin <= 24'd01045398;
                12'd2728: logsin <= 24'd01046401;
                12'd2729: logsin <= 24'd01047404;
                12'd2730: logsin <= 24'd01048409;
                12'd2731: logsin <= 24'd01049414;
                12'd2732: logsin <= 24'd01050420;
                12'd2733: logsin <= 24'd01051427;
                12'd2734: logsin <= 24'd01052434;
                12'd2735: logsin <= 24'd01053443;
                12'd2736: logsin <= 24'd01054453;
                12'd2737: logsin <= 24'd01055463;
                12'd2738: logsin <= 24'd01056475;
                12'd2739: logsin <= 24'd01057487;
                12'd2740: logsin <= 24'd01058500;
                12'd2741: logsin <= 24'd01059514;
                12'd2742: logsin <= 24'd01060529;
                12'd2743: logsin <= 24'd01061545;
                12'd2744: logsin <= 24'd01062562;
                12'd2745: logsin <= 24'd01063580;
                12'd2746: logsin <= 24'd01064598;
                12'd2747: logsin <= 24'd01065618;
                12'd2748: logsin <= 24'd01066638;
                12'd2749: logsin <= 24'd01067660;
                12'd2750: logsin <= 24'd01068682;
                12'd2751: logsin <= 24'd01069705;
                12'd2752: logsin <= 24'd01070729;
                12'd2753: logsin <= 24'd01071754;
                12'd2754: logsin <= 24'd01072780;
                12'd2755: logsin <= 24'd01073807;
                12'd2756: logsin <= 24'd01074835;
                12'd2757: logsin <= 24'd01075863;
                12'd2758: logsin <= 24'd01076893;
                12'd2759: logsin <= 24'd01077923;
                12'd2760: logsin <= 24'd01078955;
                12'd2761: logsin <= 24'd01079987;
                12'd2762: logsin <= 24'd01081021;
                12'd2763: logsin <= 24'd01082055;
                12'd2764: logsin <= 24'd01083090;
                12'd2765: logsin <= 24'd01084126;
                12'd2766: logsin <= 24'd01085163;
                12'd2767: logsin <= 24'd01086201;
                12'd2768: logsin <= 24'd01087240;
                12'd2769: logsin <= 24'd01088280;
                12'd2770: logsin <= 24'd01089321;
                12'd2771: logsin <= 24'd01090362;
                12'd2772: logsin <= 24'd01091405;
                12'd2773: logsin <= 24'd01092449;
                12'd2774: logsin <= 24'd01093493;
                12'd2775: logsin <= 24'd01094539;
                12'd2776: logsin <= 24'd01095585;
                12'd2777: logsin <= 24'd01096633;
                12'd2778: logsin <= 24'd01097681;
                12'd2779: logsin <= 24'd01098730;
                12'd2780: logsin <= 24'd01099780;
                12'd2781: logsin <= 24'd01100832;
                12'd2782: logsin <= 24'd01101884;
                12'd2783: logsin <= 24'd01102937;
                12'd2784: logsin <= 24'd01103991;
                12'd2785: logsin <= 24'd01105046;
                12'd2786: logsin <= 24'd01106102;
                12'd2787: logsin <= 24'd01107159;
                12'd2788: logsin <= 24'd01108217;
                12'd2789: logsin <= 24'd01109275;
                12'd2790: logsin <= 24'd01110335;
                12'd2791: logsin <= 24'd01111396;
                12'd2792: logsin <= 24'd01112458;
                12'd2793: logsin <= 24'd01113521;
                12'd2794: logsin <= 24'd01114584;
                12'd2795: logsin <= 24'd01115649;
                12'd2796: logsin <= 24'd01116715;
                12'd2797: logsin <= 24'd01117781;
                12'd2798: logsin <= 24'd01118849;
                12'd2799: logsin <= 24'd01119917;
                12'd2800: logsin <= 24'd01120987;
                12'd2801: logsin <= 24'd01122057;
                12'd2802: logsin <= 24'd01123129;
                12'd2803: logsin <= 24'd01124201;
                12'd2804: logsin <= 24'd01125275;
                12'd2805: logsin <= 24'd01126349;
                12'd2806: logsin <= 24'd01127425;
                12'd2807: logsin <= 24'd01128501;
                12'd2808: logsin <= 24'd01129578;
                12'd2809: logsin <= 24'd01130657;
                12'd2810: logsin <= 24'd01131736;
                12'd2811: logsin <= 24'd01132817;
                12'd2812: logsin <= 24'd01133898;
                12'd2813: logsin <= 24'd01134980;
                12'd2814: logsin <= 24'd01136064;
                12'd2815: logsin <= 24'd01137148;
                12'd2816: logsin <= 24'd01138233;
                12'd2817: logsin <= 24'd01139320;
                12'd2818: logsin <= 24'd01140407;
                12'd2819: logsin <= 24'd01141496;
                12'd2820: logsin <= 24'd01142585;
                12'd2821: logsin <= 24'd01143675;
                12'd2822: logsin <= 24'd01144767;
                12'd2823: logsin <= 24'd01145859;
                12'd2824: logsin <= 24'd01146953;
                12'd2825: logsin <= 24'd01148047;
                12'd2826: logsin <= 24'd01149142;
                12'd2827: logsin <= 24'd01150239;
                12'd2828: logsin <= 24'd01151336;
                12'd2829: logsin <= 24'd01152435;
                12'd2830: logsin <= 24'd01153534;
                12'd2831: logsin <= 24'd01154635;
                12'd2832: logsin <= 24'd01155737;
                12'd2833: logsin <= 24'd01156839;
                12'd2834: logsin <= 24'd01157943;
                12'd2835: logsin <= 24'd01159047;
                12'd2836: logsin <= 24'd01160153;
                12'd2837: logsin <= 24'd01161260;
                12'd2838: logsin <= 24'd01162368;
                12'd2839: logsin <= 24'd01163476;
                12'd2840: logsin <= 24'd01164586;
                12'd2841: logsin <= 24'd01165697;
                12'd2842: logsin <= 24'd01166809;
                12'd2843: logsin <= 24'd01167922;
                12'd2844: logsin <= 24'd01169036;
                12'd2845: logsin <= 24'd01170151;
                12'd2846: logsin <= 24'd01171267;
                12'd2847: logsin <= 24'd01172384;
                12'd2848: logsin <= 24'd01173502;
                12'd2849: logsin <= 24'd01174621;
                12'd2850: logsin <= 24'd01175742;
                12'd2851: logsin <= 24'd01176863;
                12'd2852: logsin <= 24'd01177985;
                12'd2853: logsin <= 24'd01179109;
                12'd2854: logsin <= 24'd01180233;
                12'd2855: logsin <= 24'd01181359;
                12'd2856: logsin <= 24'd01182485;
                12'd2857: logsin <= 24'd01183613;
                12'd2858: logsin <= 24'd01184742;
                12'd2859: logsin <= 24'd01185872;
                12'd2860: logsin <= 24'd01187003;
                12'd2861: logsin <= 24'd01188134;
                12'd2862: logsin <= 24'd01189267;
                12'd2863: logsin <= 24'd01190402;
                12'd2864: logsin <= 24'd01191537;
                12'd2865: logsin <= 24'd01192673;
                12'd2866: logsin <= 24'd01193810;
                12'd2867: logsin <= 24'd01194949;
                12'd2868: logsin <= 24'd01196088;
                12'd2869: logsin <= 24'd01197229;
                12'd2870: logsin <= 24'd01198370;
                12'd2871: logsin <= 24'd01199513;
                12'd2872: logsin <= 24'd01200657;
                12'd2873: logsin <= 24'd01201802;
                12'd2874: logsin <= 24'd01202948;
                12'd2875: logsin <= 24'd01204095;
                12'd2876: logsin <= 24'd01205243;
                12'd2877: logsin <= 24'd01206392;
                12'd2878: logsin <= 24'd01207542;
                12'd2879: logsin <= 24'd01208694;
                12'd2880: logsin <= 24'd01209846;
                12'd2881: logsin <= 24'd01211000;
                12'd2882: logsin <= 24'd01212155;
                12'd2883: logsin <= 24'd01213311;
                12'd2884: logsin <= 24'd01214468;
                12'd2885: logsin <= 24'd01215626;
                12'd2886: logsin <= 24'd01216785;
                12'd2887: logsin <= 24'd01217945;
                12'd2888: logsin <= 24'd01219107;
                12'd2889: logsin <= 24'd01220269;
                12'd2890: logsin <= 24'd01221433;
                12'd2891: logsin <= 24'd01222597;
                12'd2892: logsin <= 24'd01223763;
                12'd2893: logsin <= 24'd01224930;
                12'd2894: logsin <= 24'd01226098;
                12'd2895: logsin <= 24'd01227268;
                12'd2896: logsin <= 24'd01228438;
                12'd2897: logsin <= 24'd01229610;
                12'd2898: logsin <= 24'd01230782;
                12'd2899: logsin <= 24'd01231956;
                12'd2900: logsin <= 24'd01233131;
                12'd2901: logsin <= 24'd01234307;
                12'd2902: logsin <= 24'd01235484;
                12'd2903: logsin <= 24'd01236662;
                12'd2904: logsin <= 24'd01237842;
                12'd2905: logsin <= 24'd01239022;
                12'd2906: logsin <= 24'd01240204;
                12'd2907: logsin <= 24'd01241387;
                12'd2908: logsin <= 24'd01242571;
                12'd2909: logsin <= 24'd01243756;
                12'd2910: logsin <= 24'd01244943;
                12'd2911: logsin <= 24'd01246130;
                12'd2912: logsin <= 24'd01247319;
                12'd2913: logsin <= 24'd01248508;
                12'd2914: logsin <= 24'd01249699;
                12'd2915: logsin <= 24'd01250892;
                12'd2916: logsin <= 24'd01252085;
                12'd2917: logsin <= 24'd01253279;
                12'd2918: logsin <= 24'd01254475;
                12'd2919: logsin <= 24'd01255672;
                12'd2920: logsin <= 24'd01256870;
                12'd2921: logsin <= 24'd01258069;
                12'd2922: logsin <= 24'd01259269;
                12'd2923: logsin <= 24'd01260471;
                12'd2924: logsin <= 24'd01261673;
                12'd2925: logsin <= 24'd01262877;
                12'd2926: logsin <= 24'd01264082;
                12'd2927: logsin <= 24'd01265288;
                12'd2928: logsin <= 24'd01266496;
                12'd2929: logsin <= 24'd01267704;
                12'd2930: logsin <= 24'd01268914;
                12'd2931: logsin <= 24'd01270125;
                12'd2932: logsin <= 24'd01271337;
                12'd2933: logsin <= 24'd01272550;
                12'd2934: logsin <= 24'd01273765;
                12'd2935: logsin <= 24'd01274981;
                12'd2936: logsin <= 24'd01276198;
                12'd2937: logsin <= 24'd01277416;
                12'd2938: logsin <= 24'd01278635;
                12'd2939: logsin <= 24'd01279856;
                12'd2940: logsin <= 24'd01281077;
                12'd2941: logsin <= 24'd01282300;
                12'd2942: logsin <= 24'd01283525;
                12'd2943: logsin <= 24'd01284750;
                12'd2944: logsin <= 24'd01285977;
                12'd2945: logsin <= 24'd01287204;
                12'd2946: logsin <= 24'd01288433;
                12'd2947: logsin <= 24'd01289664;
                12'd2948: logsin <= 24'd01290895;
                12'd2949: logsin <= 24'd01292128;
                12'd2950: logsin <= 24'd01293362;
                12'd2951: logsin <= 24'd01294597;
                12'd2952: logsin <= 24'd01295833;
                12'd2953: logsin <= 24'd01297071;
                12'd2954: logsin <= 24'd01298310;
                12'd2955: logsin <= 24'd01299550;
                12'd2956: logsin <= 24'd01300791;
                12'd2957: logsin <= 24'd01302034;
                12'd2958: logsin <= 24'd01303278;
                12'd2959: logsin <= 24'd01304523;
                12'd2960: logsin <= 24'd01305769;
                12'd2961: logsin <= 24'd01307017;
                12'd2962: logsin <= 24'd01308266;
                12'd2963: logsin <= 24'd01309516;
                12'd2964: logsin <= 24'd01310767;
                12'd2965: logsin <= 24'd01312020;
                12'd2966: logsin <= 24'd01313274;
                12'd2967: logsin <= 24'd01314529;
                12'd2968: logsin <= 24'd01315785;
                12'd2969: logsin <= 24'd01317043;
                12'd2970: logsin <= 24'd01318302;
                12'd2971: logsin <= 24'd01319562;
                12'd2972: logsin <= 24'd01320823;
                12'd2973: logsin <= 24'd01322086;
                12'd2974: logsin <= 24'd01323350;
                12'd2975: logsin <= 24'd01324616;
                12'd2976: logsin <= 24'd01325882;
                12'd2977: logsin <= 24'd01327150;
                12'd2978: logsin <= 24'd01328419;
                12'd2979: logsin <= 24'd01329690;
                12'd2980: logsin <= 24'd01330961;
                12'd2981: logsin <= 24'd01332234;
                12'd2982: logsin <= 24'd01333509;
                12'd2983: logsin <= 24'd01334784;
                12'd2984: logsin <= 24'd01336061;
                12'd2985: logsin <= 24'd01337339;
                12'd2986: logsin <= 24'd01338619;
                12'd2987: logsin <= 24'd01339900;
                12'd2988: logsin <= 24'd01341182;
                12'd2989: logsin <= 24'd01342465;
                12'd2990: logsin <= 24'd01343750;
                12'd2991: logsin <= 24'd01345036;
                12'd2992: logsin <= 24'd01346324;
                12'd2993: logsin <= 24'd01347612;
                12'd2994: logsin <= 24'd01348902;
                12'd2995: logsin <= 24'd01350194;
                12'd2996: logsin <= 24'd01351487;
                12'd2997: logsin <= 24'd01352781;
                12'd2998: logsin <= 24'd01354076;
                12'd2999: logsin <= 24'd01355373;
                12'd3000: logsin <= 24'd01356671;
                12'd3001: logsin <= 24'd01357970;
                12'd3002: logsin <= 24'd01359271;
                12'd3003: logsin <= 24'd01360573;
                12'd3004: logsin <= 24'd01361876;
                12'd3005: logsin <= 24'd01363181;
                12'd3006: logsin <= 24'd01364487;
                12'd3007: logsin <= 24'd01365794;
                12'd3008: logsin <= 24'd01367103;
                12'd3009: logsin <= 24'd01368413;
                12'd3010: logsin <= 24'd01369725;
                12'd3011: logsin <= 24'd01371038;
                12'd3012: logsin <= 24'd01372352;
                12'd3013: logsin <= 24'd01373667;
                12'd3014: logsin <= 24'd01374984;
                12'd3015: logsin <= 24'd01376303;
                12'd3016: logsin <= 24'd01377622;
                12'd3017: logsin <= 24'd01378943;
                12'd3018: logsin <= 24'd01380266;
                12'd3019: logsin <= 24'd01381590;
                12'd3020: logsin <= 24'd01382915;
                12'd3021: logsin <= 24'd01384241;
                12'd3022: logsin <= 24'd01385569;
                12'd3023: logsin <= 24'd01386899;
                12'd3024: logsin <= 24'd01388230;
                12'd3025: logsin <= 24'd01389562;
                12'd3026: logsin <= 24'd01390895;
                12'd3027: logsin <= 24'd01392230;
                12'd3028: logsin <= 24'd01393567;
                12'd3029: logsin <= 24'd01394904;
                12'd3030: logsin <= 24'd01396243;
                12'd3031: logsin <= 24'd01397584;
                12'd3032: logsin <= 24'd01398926;
                12'd3033: logsin <= 24'd01400269;
                12'd3034: logsin <= 24'd01401614;
                12'd3035: logsin <= 24'd01402960;
                12'd3036: logsin <= 24'd01404308;
                12'd3037: logsin <= 24'd01405657;
                12'd3038: logsin <= 24'd01407008;
                12'd3039: logsin <= 24'd01408360;
                12'd3040: logsin <= 24'd01409713;
                12'd3041: logsin <= 24'd01411068;
                12'd3042: logsin <= 24'd01412424;
                12'd3043: logsin <= 24'd01413782;
                12'd3044: logsin <= 24'd01415141;
                12'd3045: logsin <= 24'd01416501;
                12'd3046: logsin <= 24'd01417863;
                12'd3047: logsin <= 24'd01419227;
                12'd3048: logsin <= 24'd01420592;
                12'd3049: logsin <= 24'd01421958;
                12'd3050: logsin <= 24'd01423326;
                12'd3051: logsin <= 24'd01424695;
                12'd3052: logsin <= 24'd01426066;
                12'd3053: logsin <= 24'd01427438;
                12'd3054: logsin <= 24'd01428812;
                12'd3055: logsin <= 24'd01430187;
                12'd3056: logsin <= 24'd01431564;
                12'd3057: logsin <= 24'd01432942;
                12'd3058: logsin <= 24'd01434322;
                12'd3059: logsin <= 24'd01435703;
                12'd3060: logsin <= 24'd01437085;
                12'd3061: logsin <= 24'd01438469;
                12'd3062: logsin <= 24'd01439855;
                12'd3063: logsin <= 24'd01441242;
                12'd3064: logsin <= 24'd01442630;
                12'd3065: logsin <= 24'd01444020;
                12'd3066: logsin <= 24'd01445412;
                12'd3067: logsin <= 24'd01446805;
                12'd3068: logsin <= 24'd01448199;
                12'd3069: logsin <= 24'd01449595;
                12'd3070: logsin <= 24'd01450993;
                12'd3071: logsin <= 24'd01452392;
                12'd3072: logsin <= 24'd01453793;
                12'd3073: logsin <= 24'd01455195;
                12'd3074: logsin <= 24'd01456598;
                12'd3075: logsin <= 24'd01458004;
                12'd3076: logsin <= 24'd01459410;
                12'd3077: logsin <= 24'd01460818;
                12'd3078: logsin <= 24'd01462228;
                12'd3079: logsin <= 24'd01463639;
                12'd3080: logsin <= 24'd01465052;
                12'd3081: logsin <= 24'd01466467;
                12'd3082: logsin <= 24'd01467883;
                12'd3083: logsin <= 24'd01469300;
                12'd3084: logsin <= 24'd01470719;
                12'd3085: logsin <= 24'd01472140;
                12'd3086: logsin <= 24'd01473562;
                12'd3087: logsin <= 24'd01474985;
                12'd3088: logsin <= 24'd01476411;
                12'd3089: logsin <= 24'd01477838;
                12'd3090: logsin <= 24'd01479266;
                12'd3091: logsin <= 24'd01480696;
                12'd3092: logsin <= 24'd01482127;
                12'd3093: logsin <= 24'd01483561;
                12'd3094: logsin <= 24'd01484995;
                12'd3095: logsin <= 24'd01486432;
                12'd3096: logsin <= 24'd01487869;
                12'd3097: logsin <= 24'd01489309;
                12'd3098: logsin <= 24'd01490750;
                12'd3099: logsin <= 24'd01492193;
                12'd3100: logsin <= 24'd01493637;
                12'd3101: logsin <= 24'd01495083;
                12'd3102: logsin <= 24'd01496530;
                12'd3103: logsin <= 24'd01497979;
                12'd3104: logsin <= 24'd01499430;
                12'd3105: logsin <= 24'd01500882;
                12'd3106: logsin <= 24'd01502336;
                12'd3107: logsin <= 24'd01503792;
                12'd3108: logsin <= 24'd01505249;
                12'd3109: logsin <= 24'd01506708;
                12'd3110: logsin <= 24'd01508168;
                12'd3111: logsin <= 24'd01509630;
                12'd3112: logsin <= 24'd01511094;
                12'd3113: logsin <= 24'd01512559;
                12'd3114: logsin <= 24'd01514026;
                12'd3115: logsin <= 24'd01515495;
                12'd3116: logsin <= 24'd01516965;
                12'd3117: logsin <= 24'd01518437;
                12'd3118: logsin <= 24'd01519911;
                12'd3119: logsin <= 24'd01521386;
                12'd3120: logsin <= 24'd01522863;
                12'd3121: logsin <= 24'd01524341;
                12'd3122: logsin <= 24'd01525822;
                12'd3123: logsin <= 24'd01527304;
                12'd3124: logsin <= 24'd01528787;
                12'd3125: logsin <= 24'd01530272;
                12'd3126: logsin <= 24'd01531759;
                12'd3127: logsin <= 24'd01533248;
                12'd3128: logsin <= 24'd01534738;
                12'd3129: logsin <= 24'd01536230;
                12'd3130: logsin <= 24'd01537724;
                12'd3131: logsin <= 24'd01539220;
                12'd3132: logsin <= 24'd01540717;
                12'd3133: logsin <= 24'd01542215;
                12'd3134: logsin <= 24'd01543716;
                12'd3135: logsin <= 24'd01545218;
                12'd3136: logsin <= 24'd01546722;
                12'd3137: logsin <= 24'd01548228;
                12'd3138: logsin <= 24'd01549735;
                12'd3139: logsin <= 24'd01551244;
                12'd3140: logsin <= 24'd01552755;
                12'd3141: logsin <= 24'd01554268;
                12'd3142: logsin <= 24'd01555782;
                12'd3143: logsin <= 24'd01557298;
                12'd3144: logsin <= 24'd01558816;
                12'd3145: logsin <= 24'd01560336;
                12'd3146: logsin <= 24'd01561857;
                12'd3147: logsin <= 24'd01563380;
                12'd3148: logsin <= 24'd01564905;
                12'd3149: logsin <= 24'd01566431;
                12'd3150: logsin <= 24'd01567960;
                12'd3151: logsin <= 24'd01569490;
                12'd3152: logsin <= 24'd01571022;
                12'd3153: logsin <= 24'd01572555;
                12'd3154: logsin <= 24'd01574091;
                12'd3155: logsin <= 24'd01575628;
                12'd3156: logsin <= 24'd01577167;
                12'd3157: logsin <= 24'd01578708;
                12'd3158: logsin <= 24'd01580251;
                12'd3159: logsin <= 24'd01581795;
                12'd3160: logsin <= 24'd01583341;
                12'd3161: logsin <= 24'd01584889;
                12'd3162: logsin <= 24'd01586439;
                12'd3163: logsin <= 24'd01587991;
                12'd3164: logsin <= 24'd01589544;
                12'd3165: logsin <= 24'd01591099;
                12'd3166: logsin <= 24'd01592656;
                12'd3167: logsin <= 24'd01594215;
                12'd3168: logsin <= 24'd01595776;
                12'd3169: logsin <= 24'd01597339;
                12'd3170: logsin <= 24'd01598903;
                12'd3171: logsin <= 24'd01600469;
                12'd3172: logsin <= 24'd01602037;
                12'd3173: logsin <= 24'd01603607;
                12'd3174: logsin <= 24'd01605179;
                12'd3175: logsin <= 24'd01606753;
                12'd3176: logsin <= 24'd01608328;
                12'd3177: logsin <= 24'd01609906;
                12'd3178: logsin <= 24'd01611485;
                12'd3179: logsin <= 24'd01613066;
                12'd3180: logsin <= 24'd01614649;
                12'd3181: logsin <= 24'd01616234;
                12'd3182: logsin <= 24'd01617821;
                12'd3183: logsin <= 24'd01619409;
                12'd3184: logsin <= 24'd01621000;
                12'd3185: logsin <= 24'd01622592;
                12'd3186: logsin <= 24'd01624187;
                12'd3187: logsin <= 24'd01625783;
                12'd3188: logsin <= 24'd01627381;
                12'd3189: logsin <= 24'd01628981;
                12'd3190: logsin <= 24'd01630583;
                12'd3191: logsin <= 24'd01632187;
                12'd3192: logsin <= 24'd01633793;
                12'd3193: logsin <= 24'd01635401;
                12'd3194: logsin <= 24'd01637010;
                12'd3195: logsin <= 24'd01638622;
                12'd3196: logsin <= 24'd01640236;
                12'd3197: logsin <= 24'd01641851;
                12'd3198: logsin <= 24'd01643469;
                12'd3199: logsin <= 24'd01645088;
                12'd3200: logsin <= 24'd01646709;
                12'd3201: logsin <= 24'd01648333;
                12'd3202: logsin <= 24'd01649958;
                12'd3203: logsin <= 24'd01651585;
                12'd3204: logsin <= 24'd01653215;
                12'd3205: logsin <= 24'd01654846;
                12'd3206: logsin <= 24'd01656479;
                12'd3207: logsin <= 24'd01658114;
                12'd3208: logsin <= 24'd01659752;
                12'd3209: logsin <= 24'd01661391;
                12'd3210: logsin <= 24'd01663032;
                12'd3211: logsin <= 24'd01664675;
                12'd3212: logsin <= 24'd01666320;
                12'd3213: logsin <= 24'd01667968;
                12'd3214: logsin <= 24'd01669617;
                12'd3215: logsin <= 24'd01671268;
                12'd3216: logsin <= 24'd01672921;
                12'd3217: logsin <= 24'd01674577;
                12'd3218: logsin <= 24'd01676234;
                12'd3219: logsin <= 24'd01677894;
                12'd3220: logsin <= 24'd01679555;
                12'd3221: logsin <= 24'd01681219;
                12'd3222: logsin <= 24'd01682884;
                12'd3223: logsin <= 24'd01684552;
                12'd3224: logsin <= 24'd01686221;
                12'd3225: logsin <= 24'd01687893;
                12'd3226: logsin <= 24'd01689567;
                12'd3227: logsin <= 24'd01691243;
                12'd3228: logsin <= 24'd01692921;
                12'd3229: logsin <= 24'd01694601;
                12'd3230: logsin <= 24'd01696283;
                12'd3231: logsin <= 24'd01697967;
                12'd3232: logsin <= 24'd01699654;
                12'd3233: logsin <= 24'd01701342;
                12'd3234: logsin <= 24'd01703033;
                12'd3235: logsin <= 24'd01704725;
                12'd3236: logsin <= 24'd01706420;
                12'd3237: logsin <= 24'd01708117;
                12'd3238: logsin <= 24'd01709816;
                12'd3239: logsin <= 24'd01711517;
                12'd3240: logsin <= 24'd01713221;
                12'd3241: logsin <= 24'd01714926;
                12'd3242: logsin <= 24'd01716634;
                12'd3243: logsin <= 24'd01718343;
                12'd3244: logsin <= 24'd01720055;
                12'd3245: logsin <= 24'd01721769;
                12'd3246: logsin <= 24'd01723486;
                12'd3247: logsin <= 24'd01725204;
                12'd3248: logsin <= 24'd01726925;
                12'd3249: logsin <= 24'd01728647;
                12'd3250: logsin <= 24'd01730372;
                12'd3251: logsin <= 24'd01732100;
                12'd3252: logsin <= 24'd01733829;
                12'd3253: logsin <= 24'd01735560;
                12'd3254: logsin <= 24'd01737294;
                12'd3255: logsin <= 24'd01739030;
                12'd3256: logsin <= 24'd01740768;
                12'd3257: logsin <= 24'd01742509;
                12'd3258: logsin <= 24'd01744251;
                12'd3259: logsin <= 24'd01745996;
                12'd3260: logsin <= 24'd01747743;
                12'd3261: logsin <= 24'd01749493;
                12'd3262: logsin <= 24'd01751244;
                12'd3263: logsin <= 24'd01752998;
                12'd3264: logsin <= 24'd01754754;
                12'd3265: logsin <= 24'd01756513;
                12'd3266: logsin <= 24'd01758273;
                12'd3267: logsin <= 24'd01760036;
                12'd3268: logsin <= 24'd01761802;
                12'd3269: logsin <= 24'd01763569;
                12'd3270: logsin <= 24'd01765339;
                12'd3271: logsin <= 24'd01767111;
                12'd3272: logsin <= 24'd01768885;
                12'd3273: logsin <= 24'd01770662;
                12'd3274: logsin <= 24'd01772441;
                12'd3275: logsin <= 24'd01774222;
                12'd3276: logsin <= 24'd01776006;
                12'd3277: logsin <= 24'd01777792;
                12'd3278: logsin <= 24'd01779580;
                12'd3279: logsin <= 24'd01781371;
                12'd3280: logsin <= 24'd01783164;
                12'd3281: logsin <= 24'd01784959;
                12'd3282: logsin <= 24'd01786757;
                12'd3283: logsin <= 24'd01788557;
                12'd3284: logsin <= 24'd01790359;
                12'd3285: logsin <= 24'd01792164;
                12'd3286: logsin <= 24'd01793971;
                12'd3287: logsin <= 24'd01795781;
                12'd3288: logsin <= 24'd01797593;
                12'd3289: logsin <= 24'd01799407;
                12'd3290: logsin <= 24'd01801224;
                12'd3291: logsin <= 24'd01803043;
                12'd3292: logsin <= 24'd01804864;
                12'd3293: logsin <= 24'd01806688;
                12'd3294: logsin <= 24'd01808515;
                12'd3295: logsin <= 24'd01810344;
                12'd3296: logsin <= 24'd01812175;
                12'd3297: logsin <= 24'd01814009;
                12'd3298: logsin <= 24'd01815845;
                12'd3299: logsin <= 24'd01817683;
                12'd3300: logsin <= 24'd01819524;
                12'd3301: logsin <= 24'd01821368;
                12'd3302: logsin <= 24'd01823214;
                12'd3303: logsin <= 24'd01825062;
                12'd3304: logsin <= 24'd01826913;
                12'd3305: logsin <= 24'd01828767;
                12'd3306: logsin <= 24'd01830623;
                12'd3307: logsin <= 24'd01832481;
                12'd3308: logsin <= 24'd01834342;
                12'd3309: logsin <= 24'd01836206;
                12'd3310: logsin <= 24'd01838072;
                12'd3311: logsin <= 24'd01839940;
                12'd3312: logsin <= 24'd01841811;
                12'd3313: logsin <= 24'd01843685;
                12'd3314: logsin <= 24'd01845561;
                12'd3315: logsin <= 24'd01847440;
                12'd3316: logsin <= 24'd01849321;
                12'd3317: logsin <= 24'd01851205;
                12'd3318: logsin <= 24'd01853091;
                12'd3319: logsin <= 24'd01854980;
                12'd3320: logsin <= 24'd01856872;
                12'd3321: logsin <= 24'd01858766;
                12'd3322: logsin <= 24'd01860663;
                12'd3323: logsin <= 24'd01862562;
                12'd3324: logsin <= 24'd01864464;
                12'd3325: logsin <= 24'd01866369;
                12'd3326: logsin <= 24'd01868276;
                12'd3327: logsin <= 24'd01870186;
                12'd3328: logsin <= 24'd01872098;
                12'd3329: logsin <= 24'd01874013;
                12'd3330: logsin <= 24'd01875931;
                12'd3331: logsin <= 24'd01877851;
                12'd3332: logsin <= 24'd01879775;
                12'd3333: logsin <= 24'd01881700;
                12'd3334: logsin <= 24'd01883629;
                12'd3335: logsin <= 24'd01885560;
                12'd3336: logsin <= 24'd01887494;
                12'd3337: logsin <= 24'd01889430;
                12'd3338: logsin <= 24'd01891369;
                12'd3339: logsin <= 24'd01893311;
                12'd3340: logsin <= 24'd01895256;
                12'd3341: logsin <= 24'd01897203;
                12'd3342: logsin <= 24'd01899153;
                12'd3343: logsin <= 24'd01901106;
                12'd3344: logsin <= 24'd01903062;
                12'd3345: logsin <= 24'd01905020;
                12'd3346: logsin <= 24'd01906981;
                12'd3347: logsin <= 24'd01908945;
                12'd3348: logsin <= 24'd01910912;
                12'd3349: logsin <= 24'd01912881;
                12'd3350: logsin <= 24'd01914853;
                12'd3351: logsin <= 24'd01916829;
                12'd3352: logsin <= 24'd01918806;
                12'd3353: logsin <= 24'd01920787;
                12'd3354: logsin <= 24'd01922770;
                12'd3355: logsin <= 24'd01924757;
                12'd3356: logsin <= 24'd01926746;
                12'd3357: logsin <= 24'd01928738;
                12'd3358: logsin <= 24'd01930733;
                12'd3359: logsin <= 24'd01932730;
                12'd3360: logsin <= 24'd01934731;
                12'd3361: logsin <= 24'd01936734;
                12'd3362: logsin <= 24'd01938740;
                12'd3363: logsin <= 24'd01940750;
                12'd3364: logsin <= 24'd01942762;
                12'd3365: logsin <= 24'd01944777;
                12'd3366: logsin <= 24'd01946795;
                12'd3367: logsin <= 24'd01948815;
                12'd3368: logsin <= 24'd01950839;
                12'd3369: logsin <= 24'd01952866;
                12'd3370: logsin <= 24'd01954895;
                12'd3371: logsin <= 24'd01956928;
                12'd3372: logsin <= 24'd01958963;
                12'd3373: logsin <= 24'd01961002;
                12'd3374: logsin <= 24'd01963043;
                12'd3375: logsin <= 24'd01965088;
                12'd3376: logsin <= 24'd01967135;
                12'd3377: logsin <= 24'd01969185;
                12'd3378: logsin <= 24'd01971239;
                12'd3379: logsin <= 24'd01973295;
                12'd3380: logsin <= 24'd01975355;
                12'd3381: logsin <= 24'd01977417;
                12'd3382: logsin <= 24'd01979483;
                12'd3383: logsin <= 24'd01981551;
                12'd3384: logsin <= 24'd01983623;
                12'd3385: logsin <= 24'd01985698;
                12'd3386: logsin <= 24'd01987775;
                12'd3387: logsin <= 24'd01989856;
                12'd3388: logsin <= 24'd01991940;
                12'd3389: logsin <= 24'd01994027;
                12'd3390: logsin <= 24'd01996117;
                12'd3391: logsin <= 24'd01998210;
                12'd3392: logsin <= 24'd02000307;
                12'd3393: logsin <= 24'd02002406;
                12'd3394: logsin <= 24'd02004509;
                12'd3395: logsin <= 24'd02006615;
                12'd3396: logsin <= 24'd02008724;
                12'd3397: logsin <= 24'd02010836;
                12'd3398: logsin <= 24'd02012951;
                12'd3399: logsin <= 24'd02015070;
                12'd3400: logsin <= 24'd02017191;
                12'd3401: logsin <= 24'd02019316;
                12'd3402: logsin <= 24'd02021444;
                12'd3403: logsin <= 24'd02023575;
                12'd3404: logsin <= 24'd02025710;
                12'd3405: logsin <= 24'd02027848;
                12'd3406: logsin <= 24'd02029989;
                12'd3407: logsin <= 24'd02032133;
                12'd3408: logsin <= 24'd02034281;
                12'd3409: logsin <= 24'd02036431;
                12'd3410: logsin <= 24'd02038586;
                12'd3411: logsin <= 24'd02040743;
                12'd3412: logsin <= 24'd02042904;
                12'd3413: logsin <= 24'd02045068;
                12'd3414: logsin <= 24'd02047235;
                12'd3415: logsin <= 24'd02049406;
                12'd3416: logsin <= 24'd02051580;
                12'd3417: logsin <= 24'd02053757;
                12'd3418: logsin <= 24'd02055938;
                12'd3419: logsin <= 24'd02058122;
                12'd3420: logsin <= 24'd02060309;
                12'd3421: logsin <= 24'd02062500;
                12'd3422: logsin <= 24'd02064694;
                12'd3423: logsin <= 24'd02066892;
                12'd3424: logsin <= 24'd02069093;
                12'd3425: logsin <= 24'd02071298;
                12'd3426: logsin <= 24'd02073506;
                12'd3427: logsin <= 24'd02075717;
                12'd3428: logsin <= 24'd02077932;
                12'd3429: logsin <= 24'd02080150;
                12'd3430: logsin <= 24'd02082372;
                12'd3431: logsin <= 24'd02084598;
                12'd3432: logsin <= 24'd02086826;
                12'd3433: logsin <= 24'd02089059;
                12'd3434: logsin <= 24'd02091295;
                12'd3435: logsin <= 24'd02093534;
                12'd3436: logsin <= 24'd02095777;
                12'd3437: logsin <= 24'd02098023;
                12'd3438: logsin <= 24'd02100273;
                12'd3439: logsin <= 24'd02102527;
                12'd3440: logsin <= 24'd02104784;
                12'd3441: logsin <= 24'd02107045;
                12'd3442: logsin <= 24'd02109309;
                12'd3443: logsin <= 24'd02111577;
                12'd3444: logsin <= 24'd02113849;
                12'd3445: logsin <= 24'd02116124;
                12'd3446: logsin <= 24'd02118403;
                12'd3447: logsin <= 24'd02120686;
                12'd3448: logsin <= 24'd02122972;
                12'd3449: logsin <= 24'd02125262;
                12'd3450: logsin <= 24'd02127556;
                12'd3451: logsin <= 24'd02129853;
                12'd3452: logsin <= 24'd02132154;
                12'd3453: logsin <= 24'd02134459;
                12'd3454: logsin <= 24'd02136768;
                12'd3455: logsin <= 24'd02139080;
                12'd3456: logsin <= 24'd02141396;
                12'd3457: logsin <= 24'd02143716;
                12'd3458: logsin <= 24'd02146039;
                12'd3459: logsin <= 24'd02148367;
                12'd3460: logsin <= 24'd02150698;
                12'd3461: logsin <= 24'd02153033;
                12'd3462: logsin <= 24'd02155372;
                12'd3463: logsin <= 24'd02157715;
                12'd3464: logsin <= 24'd02160061;
                12'd3465: logsin <= 24'd02162412;
                12'd3466: logsin <= 24'd02164766;
                12'd3467: logsin <= 24'd02167124;
                12'd3468: logsin <= 24'd02169486;
                12'd3469: logsin <= 24'd02171852;
                12'd3470: logsin <= 24'd02174222;
                12'd3471: logsin <= 24'd02176596;
                12'd3472: logsin <= 24'd02178974;
                12'd3473: logsin <= 24'd02181356;
                12'd3474: logsin <= 24'd02183742;
                12'd3475: logsin <= 24'd02186132;
                12'd3476: logsin <= 24'd02188525;
                12'd3477: logsin <= 24'd02190923;
                12'd3478: logsin <= 24'd02193325;
                12'd3479: logsin <= 24'd02195731;
                12'd3480: logsin <= 24'd02198141;
                12'd3481: logsin <= 24'd02200555;
                12'd3482: logsin <= 24'd02202973;
                12'd3483: logsin <= 24'd02205395;
                12'd3484: logsin <= 24'd02207822;
                12'd3485: logsin <= 24'd02210252;
                12'd3486: logsin <= 24'd02212687;
                12'd3487: logsin <= 24'd02215125;
                12'd3488: logsin <= 24'd02217568;
                12'd3489: logsin <= 24'd02220015;
                12'd3490: logsin <= 24'd02222466;
                12'd3491: logsin <= 24'd02224922;
                12'd3492: logsin <= 24'd02227381;
                12'd3493: logsin <= 24'd02229845;
                12'd3494: logsin <= 24'd02232313;
                12'd3495: logsin <= 24'd02234786;
                12'd3496: logsin <= 24'd02237262;
                12'd3497: logsin <= 24'd02239743;
                12'd3498: logsin <= 24'd02242229;
                12'd3499: logsin <= 24'd02244718;
                12'd3500: logsin <= 24'd02247212;
                12'd3501: logsin <= 24'd02249710;
                12'd3502: logsin <= 24'd02252213;
                12'd3503: logsin <= 24'd02254720;
                12'd3504: logsin <= 24'd02257231;
                12'd3505: logsin <= 24'd02259747;
                12'd3506: logsin <= 24'd02262267;
                12'd3507: logsin <= 24'd02264791;
                12'd3508: logsin <= 24'd02267320;
                12'd3509: logsin <= 24'd02269854;
                12'd3510: logsin <= 24'd02272392;
                12'd3511: logsin <= 24'd02274934;
                12'd3512: logsin <= 24'd02277481;
                12'd3513: logsin <= 24'd02280032;
                12'd3514: logsin <= 24'd02282588;
                12'd3515: logsin <= 24'd02285149;
                12'd3516: logsin <= 24'd02287714;
                12'd3517: logsin <= 24'd02290284;
                12'd3518: logsin <= 24'd02292858;
                12'd3519: logsin <= 24'd02295437;
                12'd3520: logsin <= 24'd02298020;
                12'd3521: logsin <= 24'd02300608;
                12'd3522: logsin <= 24'd02303201;
                12'd3523: logsin <= 24'd02305799;
                12'd3524: logsin <= 24'd02308401;
                12'd3525: logsin <= 24'd02311008;
                12'd3526: logsin <= 24'd02313619;
                12'd3527: logsin <= 24'd02316236;
                12'd3528: logsin <= 24'd02318857;
                12'd3529: logsin <= 24'd02321483;
                12'd3530: logsin <= 24'd02324113;
                12'd3531: logsin <= 24'd02326749;
                12'd3532: logsin <= 24'd02329389;
                12'd3533: logsin <= 24'd02332034;
                12'd3534: logsin <= 24'd02334684;
                12'd3535: logsin <= 24'd02337339;
                12'd3536: logsin <= 24'd02339999;
                12'd3537: logsin <= 24'd02342663;
                12'd3538: logsin <= 24'd02345333;
                12'd3539: logsin <= 24'd02348007;
                12'd3540: logsin <= 24'd02350687;
                12'd3541: logsin <= 24'd02353371;
                12'd3542: logsin <= 24'd02356061;
                12'd3543: logsin <= 24'd02358755;
                12'd3544: logsin <= 24'd02361454;
                12'd3545: logsin <= 24'd02364159;
                12'd3546: logsin <= 24'd02366869;
                12'd3547: logsin <= 24'd02369583;
                12'd3548: logsin <= 24'd02372303;
                12'd3549: logsin <= 24'd02375028;
                12'd3550: logsin <= 24'd02377758;
                12'd3551: logsin <= 24'd02380493;
                12'd3552: logsin <= 24'd02383234;
                12'd3553: logsin <= 24'd02385979;
                12'd3554: logsin <= 24'd02388730;
                12'd3555: logsin <= 24'd02391486;
                12'd3556: logsin <= 24'd02394247;
                12'd3557: logsin <= 24'd02397014;
                12'd3558: logsin <= 24'd02399786;
                12'd3559: logsin <= 24'd02402563;
                12'd3560: logsin <= 24'd02405345;
                12'd3561: logsin <= 24'd02408133;
                12'd3562: logsin <= 24'd02410926;
                12'd3563: logsin <= 24'd02413725;
                12'd3564: logsin <= 24'd02416529;
                12'd3565: logsin <= 24'd02419338;
                12'd3566: logsin <= 24'd02422153;
                12'd3567: logsin <= 24'd02424974;
                12'd3568: logsin <= 24'd02427799;
                12'd3569: logsin <= 24'd02430631;
                12'd3570: logsin <= 24'd02433468;
                12'd3571: logsin <= 24'd02436310;
                12'd3572: logsin <= 24'd02439158;
                12'd3573: logsin <= 24'd02442012;
                12'd3574: logsin <= 24'd02444871;
                12'd3575: logsin <= 24'd02447736;
                12'd3576: logsin <= 24'd02450606;
                12'd3577: logsin <= 24'd02453482;
                12'd3578: logsin <= 24'd02456364;
                12'd3579: logsin <= 24'd02459252;
                12'd3580: logsin <= 24'd02462145;
                12'd3581: logsin <= 24'd02465044;
                12'd3582: logsin <= 24'd02467949;
                12'd3583: logsin <= 24'd02470860;
                12'd3584: logsin <= 24'd02473777;
                12'd3585: logsin <= 24'd02476699;
                12'd3586: logsin <= 24'd02479627;
                12'd3587: logsin <= 24'd02482562;
                12'd3588: logsin <= 24'd02485502;
                12'd3589: logsin <= 24'd02488448;
                12'd3590: logsin <= 24'd02491400;
                12'd3591: logsin <= 24'd02494358;
                12'd3592: logsin <= 24'd02497322;
                12'd3593: logsin <= 24'd02500292;
                12'd3594: logsin <= 24'd02503268;
                12'd3595: logsin <= 24'd02506251;
                12'd3596: logsin <= 24'd02509239;
                12'd3597: logsin <= 24'd02512234;
                12'd3598: logsin <= 24'd02515234;
                12'd3599: logsin <= 24'd02518241;
                12'd3600: logsin <= 24'd02521254;
                12'd3601: logsin <= 24'd02524273;
                12'd3602: logsin <= 24'd02527299;
                12'd3603: logsin <= 24'd02530331;
                12'd3604: logsin <= 24'd02533369;
                12'd3605: logsin <= 24'd02536414;
                12'd3606: logsin <= 24'd02539464;
                12'd3607: logsin <= 24'd02542522;
                12'd3608: logsin <= 24'd02545585;
                12'd3609: logsin <= 24'd02548655;
                12'd3610: logsin <= 24'd02551732;
                12'd3611: logsin <= 24'd02554815;
                12'd3612: logsin <= 24'd02557905;
                12'd3613: logsin <= 24'd02561001;
                12'd3614: logsin <= 24'd02564104;
                12'd3615: logsin <= 24'd02567213;
                12'd3616: logsin <= 24'd02570329;
                12'd3617: logsin <= 24'd02573451;
                12'd3618: logsin <= 24'd02576581;
                12'd3619: logsin <= 24'd02579717;
                12'd3620: logsin <= 24'd02582859;
                12'd3621: logsin <= 24'd02586009;
                12'd3622: logsin <= 24'd02589165;
                12'd3623: logsin <= 24'd02592328;
                12'd3624: logsin <= 24'd02595498;
                12'd3625: logsin <= 24'd02598675;
                12'd3626: logsin <= 24'd02601859;
                12'd3627: logsin <= 24'd02605049;
                12'd3628: logsin <= 24'd02608247;
                12'd3629: logsin <= 24'd02611452;
                12'd3630: logsin <= 24'd02614663;
                12'd3631: logsin <= 24'd02617882;
                12'd3632: logsin <= 24'd02621108;
                12'd3633: logsin <= 24'd02624341;
                12'd3634: logsin <= 24'd02627581;
                12'd3635: logsin <= 24'd02630828;
                12'd3636: logsin <= 24'd02634083;
                12'd3637: logsin <= 24'd02637344;
                12'd3638: logsin <= 24'd02640613;
                12'd3639: logsin <= 24'd02643890;
                12'd3640: logsin <= 24'd02647173;
                12'd3641: logsin <= 24'd02650464;
                12'd3642: logsin <= 24'd02653763;
                12'd3643: logsin <= 24'd02657068;
                12'd3644: logsin <= 24'd02660382;
                12'd3645: logsin <= 24'd02663702;
                12'd3646: logsin <= 24'd02667031;
                12'd3647: logsin <= 24'd02670367;
                12'd3648: logsin <= 24'd02673710;
                12'd3649: logsin <= 24'd02677061;
                12'd3650: logsin <= 24'd02680420;
                12'd3651: logsin <= 24'd02683786;
                12'd3652: logsin <= 24'd02687160;
                12'd3653: logsin <= 24'd02690542;
                12'd3654: logsin <= 24'd02693932;
                12'd3655: logsin <= 24'd02697330;
                12'd3656: logsin <= 24'd02700735;
                12'd3657: logsin <= 24'd02704148;
                12'd3658: logsin <= 24'd02707570;
                12'd3659: logsin <= 24'd02710999;
                12'd3660: logsin <= 24'd02714436;
                12'd3661: logsin <= 24'd02717882;
                12'd3662: logsin <= 24'd02721335;
                12'd3663: logsin <= 24'd02724796;
                12'd3664: logsin <= 24'd02728266;
                12'd3665: logsin <= 24'd02731744;
                12'd3666: logsin <= 24'd02735230;
                12'd3667: logsin <= 24'd02738725;
                12'd3668: logsin <= 24'd02742227;
                12'd3669: logsin <= 24'd02745738;
                12'd3670: logsin <= 24'd02749258;
                12'd3671: logsin <= 24'd02752786;
                12'd3672: logsin <= 24'd02756322;
                12'd3673: logsin <= 24'd02759867;
                12'd3674: logsin <= 24'd02763420;
                12'd3675: logsin <= 24'd02766982;
                12'd3676: logsin <= 24'd02770553;
                12'd3677: logsin <= 24'd02774132;
                12'd3678: logsin <= 24'd02777720;
                12'd3679: logsin <= 24'd02781317;
                12'd3680: logsin <= 24'd02784923;
                12'd3681: logsin <= 24'd02788537;
                12'd3682: logsin <= 24'd02792161;
                12'd3683: logsin <= 24'd02795793;
                12'd3684: logsin <= 24'd02799434;
                12'd3685: logsin <= 24'd02803084;
                12'd3686: logsin <= 24'd02806743;
                12'd3687: logsin <= 24'd02810412;
                12'd3688: logsin <= 24'd02814089;
                12'd3689: logsin <= 24'd02817776;
                12'd3690: logsin <= 24'd02821472;
                12'd3691: logsin <= 24'd02825177;
                12'd3692: logsin <= 24'd02828891;
                12'd3693: logsin <= 24'd02832615;
                12'd3694: logsin <= 24'd02836349;
                12'd3695: logsin <= 24'd02840091;
                12'd3696: logsin <= 24'd02843843;
                12'd3697: logsin <= 24'd02847605;
                12'd3698: logsin <= 24'd02851377;
                12'd3699: logsin <= 24'd02855158;
                12'd3700: logsin <= 24'd02858948;
                12'd3701: logsin <= 24'd02862749;
                12'd3702: logsin <= 24'd02866559;
                12'd3703: logsin <= 24'd02870379;
                12'd3704: logsin <= 24'd02874209;
                12'd3705: logsin <= 24'd02878049;
                12'd3706: logsin <= 24'd02881899;
                12'd3707: logsin <= 24'd02885759;
                12'd3708: logsin <= 24'd02889629;
                12'd3709: logsin <= 24'd02893509;
                12'd3710: logsin <= 24'd02897400;
                12'd3711: logsin <= 24'd02901301;
                12'd3712: logsin <= 24'd02905212;
                12'd3713: logsin <= 24'd02909133;
                12'd3714: logsin <= 24'd02913065;
                12'd3715: logsin <= 24'd02917007;
                12'd3716: logsin <= 24'd02920960;
                12'd3717: logsin <= 24'd02924923;
                12'd3718: logsin <= 24'd02928897;
                12'd3719: logsin <= 24'd02932882;
                12'd3720: logsin <= 24'd02936877;
                12'd3721: logsin <= 24'd02940883;
                12'd3722: logsin <= 24'd02944900;
                12'd3723: logsin <= 24'd02948928;
                12'd3724: logsin <= 24'd02952967;
                12'd3725: logsin <= 24'd02957017;
                12'd3726: logsin <= 24'd02961079;
                12'd3727: logsin <= 24'd02965151;
                12'd3728: logsin <= 24'd02969234;
                12'd3729: logsin <= 24'd02973329;
                12'd3730: logsin <= 24'd02977435;
                12'd3731: logsin <= 24'd02981553;
                12'd3732: logsin <= 24'd02985682;
                12'd3733: logsin <= 24'd02989822;
                12'd3734: logsin <= 24'd02993974;
                12'd3735: logsin <= 24'd02998138;
                12'd3736: logsin <= 24'd03002313;
                12'd3737: logsin <= 24'd03006500;
                12'd3738: logsin <= 24'd03010700;
                12'd3739: logsin <= 24'd03014910;
                12'd3740: logsin <= 24'd03019133;
                12'd3741: logsin <= 24'd03023368;
                12'd3742: logsin <= 24'd03027616;
                12'd3743: logsin <= 24'd03031875;
                12'd3744: logsin <= 24'd03036146;
                12'd3745: logsin <= 24'd03040430;
                12'd3746: logsin <= 24'd03044726;
                12'd3747: logsin <= 24'd03049035;
                12'd3748: logsin <= 24'd03053356;
                12'd3749: logsin <= 24'd03057690;
                12'd3750: logsin <= 24'd03062037;
                12'd3751: logsin <= 24'd03066396;
                12'd3752: logsin <= 24'd03070768;
                12'd3753: logsin <= 24'd03075153;
                12'd3754: logsin <= 24'd03079551;
                12'd3755: logsin <= 24'd03083962;
                12'd3756: logsin <= 24'd03088386;
                12'd3757: logsin <= 24'd03092823;
                12'd3758: logsin <= 24'd03097274;
                12'd3759: logsin <= 24'd03101738;
                12'd3760: logsin <= 24'd03106215;
                12'd3761: logsin <= 24'd03110706;
                12'd3762: logsin <= 24'd03115210;
                12'd3763: logsin <= 24'd03119729;
                12'd3764: logsin <= 24'd03124260;
                12'd3765: logsin <= 24'd03128806;
                12'd3766: logsin <= 24'd03133366;
                12'd3767: logsin <= 24'd03137940;
                12'd3768: logsin <= 24'd03142527;
                12'd3769: logsin <= 24'd03147129;
                12'd3770: logsin <= 24'd03151746;
                12'd3771: logsin <= 24'd03156376;
                12'd3772: logsin <= 24'd03161021;
                12'd3773: logsin <= 24'd03165681;
                12'd3774: logsin <= 24'd03170355;
                12'd3775: logsin <= 24'd03175044;
                12'd3776: logsin <= 24'd03179747;
                12'd3777: logsin <= 24'd03184466;
                12'd3778: logsin <= 24'd03189199;
                12'd3779: logsin <= 24'd03193948;
                12'd3780: logsin <= 24'd03198712;
                12'd3781: logsin <= 24'd03203491;
                12'd3782: logsin <= 24'd03208285;
                12'd3783: logsin <= 24'd03213095;
                12'd3784: logsin <= 24'd03217921;
                12'd3785: logsin <= 24'd03222762;
                12'd3786: logsin <= 24'd03227619;
                12'd3787: logsin <= 24'd03232492;
                12'd3788: logsin <= 24'd03237380;
                12'd3789: logsin <= 24'd03242285;
                12'd3790: logsin <= 24'd03247206;
                12'd3791: logsin <= 24'd03252144;
                12'd3792: logsin <= 24'd03257097;
                12'd3793: logsin <= 24'd03262067;
                12'd3794: logsin <= 24'd03267054;
                12'd3795: logsin <= 24'd03272058;
                12'd3796: logsin <= 24'd03277078;
                12'd3797: logsin <= 24'd03282115;
                12'd3798: logsin <= 24'd03287170;
                12'd3799: logsin <= 24'd03292241;
                12'd3800: logsin <= 24'd03297330;
                12'd3801: logsin <= 24'd03302436;
                12'd3802: logsin <= 24'd03307560;
                12'd3803: logsin <= 24'd03312701;
                12'd3804: logsin <= 24'd03317860;
                12'd3805: logsin <= 24'd03323037;
                12'd3806: logsin <= 24'd03328232;
                12'd3807: logsin <= 24'd03333445;
                12'd3808: logsin <= 24'd03338676;
                12'd3809: logsin <= 24'd03343926;
                12'd3810: logsin <= 24'd03349194;
                12'd3811: logsin <= 24'd03354481;
                12'd3812: logsin <= 24'd03359787;
                12'd3813: logsin <= 24'd03365111;
                12'd3814: logsin <= 24'd03370455;
                12'd3815: logsin <= 24'd03375817;
                12'd3816: logsin <= 24'd03381199;
                12'd3817: logsin <= 24'd03386601;
                12'd3818: logsin <= 24'd03392022;
                12'd3819: logsin <= 24'd03397463;
                12'd3820: logsin <= 24'd03402923;
                12'd3821: logsin <= 24'd03408404;
                12'd3822: logsin <= 24'd03413904;
                12'd3823: logsin <= 24'd03419426;
                12'd3824: logsin <= 24'd03424967;
                12'd3825: logsin <= 24'd03430529;
                12'd3826: logsin <= 24'd03436112;
                12'd3827: logsin <= 24'd03441716;
                12'd3828: logsin <= 24'd03447340;
                12'd3829: logsin <= 24'd03452987;
                12'd3830: logsin <= 24'd03458654;
                12'd3831: logsin <= 24'd03464343;
                12'd3832: logsin <= 24'd03470053;
                12'd3833: logsin <= 24'd03475786;
                12'd3834: logsin <= 24'd03481540;
                12'd3835: logsin <= 24'd03487317;
                12'd3836: logsin <= 24'd03493116;
                12'd3837: logsin <= 24'd03498938;
                12'd3838: logsin <= 24'd03504782;
                12'd3839: logsin <= 24'd03510649;
                12'd3840: logsin <= 24'd03516540;
                12'd3841: logsin <= 24'd03522453;
                12'd3842: logsin <= 24'd03528390;
                12'd3843: logsin <= 24'd03534351;
                12'd3844: logsin <= 24'd03540335;
                12'd3845: logsin <= 24'd03546344;
                12'd3846: logsin <= 24'd03552376;
                12'd3847: logsin <= 24'd03558433;
                12'd3848: logsin <= 24'd03564515;
                12'd3849: logsin <= 24'd03570621;
                12'd3850: logsin <= 24'd03576752;
                12'd3851: logsin <= 24'd03582909;
                12'd3852: logsin <= 24'd03589090;
                12'd3853: logsin <= 24'd03595298;
                12'd3854: logsin <= 24'd03601531;
                12'd3855: logsin <= 24'd03607790;
                12'd3856: logsin <= 24'd03614076;
                12'd3857: logsin <= 24'd03620387;
                12'd3858: logsin <= 24'd03626726;
                12'd3859: logsin <= 24'd03633091;
                12'd3860: logsin <= 24'd03639484;
                12'd3861: logsin <= 24'd03645904;
                12'd3862: logsin <= 24'd03652351;
                12'd3863: logsin <= 24'd03658827;
                12'd3864: logsin <= 24'd03665330;
                12'd3865: logsin <= 24'd03671862;
                12'd3866: logsin <= 24'd03678422;
                12'd3867: logsin <= 24'd03685011;
                12'd3868: logsin <= 24'd03691629;
                12'd3869: logsin <= 24'd03698276;
                12'd3870: logsin <= 24'd03704953;
                12'd3871: logsin <= 24'd03711660;
                12'd3872: logsin <= 24'd03718397;
                12'd3873: logsin <= 24'd03725164;
                12'd3874: logsin <= 24'd03731962;
                12'd3875: logsin <= 24'd03738791;
                12'd3876: logsin <= 24'd03745651;
                12'd3877: logsin <= 24'd03752542;
                12'd3878: logsin <= 24'd03759465;
                12'd3879: logsin <= 24'd03766421;
                12'd3880: logsin <= 24'd03773408;
                12'd3881: logsin <= 24'd03780428;
                12'd3882: logsin <= 24'd03787482;
                12'd3883: logsin <= 24'd03794568;
                12'd3884: logsin <= 24'd03801688;
                12'd3885: logsin <= 24'd03808842;
                12'd3886: logsin <= 24'd03816030;
                12'd3887: logsin <= 24'd03823253;
                12'd3888: logsin <= 24'd03830510;
                12'd3889: logsin <= 24'd03837803;
                12'd3890: logsin <= 24'd03845131;
                12'd3891: logsin <= 24'd03852495;
                12'd3892: logsin <= 24'd03859896;
                12'd3893: logsin <= 24'd03867333;
                12'd3894: logsin <= 24'd03874807;
                12'd3895: logsin <= 24'd03882318;
                12'd3896: logsin <= 24'd03889867;
                12'd3897: logsin <= 24'd03897455;
                12'd3898: logsin <= 24'd03905080;
                12'd3899: logsin <= 24'd03912745;
                12'd3900: logsin <= 24'd03920448;
                12'd3901: logsin <= 24'd03928192;
                12'd3902: logsin <= 24'd03935975;
                12'd3903: logsin <= 24'd03943799;
                12'd3904: logsin <= 24'd03951664;
                12'd3905: logsin <= 24'd03959570;
                12'd3906: logsin <= 24'd03967518;
                12'd3907: logsin <= 24'd03975508;
                12'd3908: logsin <= 24'd03983541;
                12'd3909: logsin <= 24'd03991617;
                12'd3910: logsin <= 24'd03999736;
                12'd3911: logsin <= 24'd04007899;
                12'd3912: logsin <= 24'd04016107;
                12'd3913: logsin <= 24'd04024360;
                12'd3914: logsin <= 24'd04032659;
                12'd3915: logsin <= 24'd04041003;
                12'd3916: logsin <= 24'd04049394;
                12'd3917: logsin <= 24'd04057832;
                12'd3918: logsin <= 24'd04066318;
                12'd3919: logsin <= 24'd04074852;
                12'd3920: logsin <= 24'd04083434;
                12'd3921: logsin <= 24'd04092065;
                12'd3922: logsin <= 24'd04100747;
                12'd3923: logsin <= 24'd04109478;
                12'd3924: logsin <= 24'd04118261;
                12'd3925: logsin <= 24'd04127095;
                12'd3926: logsin <= 24'd04135981;
                12'd3927: logsin <= 24'd04144919;
                12'd3928: logsin <= 24'd04153912;
                12'd3929: logsin <= 24'd04162958;
                12'd3930: logsin <= 24'd04172059;
                12'd3931: logsin <= 24'd04181215;
                12'd3932: logsin <= 24'd04190427;
                12'd3933: logsin <= 24'd04199696;
                12'd3934: logsin <= 24'd04209022;
                12'd3935: logsin <= 24'd04218406;
                12'd3936: logsin <= 24'd04227849;
                12'd3937: logsin <= 24'd04237352;
                12'd3938: logsin <= 24'd04246914;
                12'd3939: logsin <= 24'd04256538;
                12'd3940: logsin <= 24'd04266224;
                12'd3941: logsin <= 24'd04275972;
                12'd3942: logsin <= 24'd04285784;
                12'd3943: logsin <= 24'd04295660;
                12'd3944: logsin <= 24'd04305602;
                12'd3945: logsin <= 24'd04315609;
                12'd3946: logsin <= 24'd04325683;
                12'd3947: logsin <= 24'd04335825;
                12'd3948: logsin <= 24'd04346035;
                12'd3949: logsin <= 24'd04356315;
                12'd3950: logsin <= 24'd04366666;
                12'd3951: logsin <= 24'd04377088;
                12'd3952: logsin <= 24'd04387583;
                12'd3953: logsin <= 24'd04398151;
                12'd3954: logsin <= 24'd04408794;
                12'd3955: logsin <= 24'd04419513;
                12'd3956: logsin <= 24'd04430308;
                12'd3957: logsin <= 24'd04441181;
                12'd3958: logsin <= 24'd04452133;
                12'd3959: logsin <= 24'd04463165;
                12'd3960: logsin <= 24'd04474278;
                12'd3961: logsin <= 24'd04485474;
                12'd3962: logsin <= 24'd04496753;
                12'd3963: logsin <= 24'd04508118;
                12'd3964: logsin <= 24'd04519569;
                12'd3965: logsin <= 24'd04531107;
                12'd3966: logsin <= 24'd04542734;
                12'd3967: logsin <= 24'd04554451;
                12'd3968: logsin <= 24'd04566260;
                12'd3969: logsin <= 24'd04578163;
                12'd3970: logsin <= 24'd04590160;
                12'd3971: logsin <= 24'd04602253;
                12'd3972: logsin <= 24'd04614443;
                12'd3973: logsin <= 24'd04626733;
                12'd3974: logsin <= 24'd04639124;
                12'd3975: logsin <= 24'd04651617;
                12'd3976: logsin <= 24'd04664215;
                12'd3977: logsin <= 24'd04676919;
                12'd3978: logsin <= 24'd04689730;
                12'd3979: logsin <= 24'd04702651;
                12'd3980: logsin <= 24'd04715684;
                12'd3981: logsin <= 24'd04728830;
                12'd3982: logsin <= 24'd04742092;
                12'd3983: logsin <= 24'd04755471;
                12'd3984: logsin <= 24'd04768969;
                12'd3985: logsin <= 24'd04782590;
                12'd3986: logsin <= 24'd04796334;
                12'd3987: logsin <= 24'd04810205;
                12'd3988: logsin <= 24'd04824204;
                12'd3989: logsin <= 24'd04838335;
                12'd3990: logsin <= 24'd04852598;
                12'd3991: logsin <= 24'd04866998;
                12'd3992: logsin <= 24'd04881536;
                12'd3993: logsin <= 24'd04896216;
                12'd3994: logsin <= 24'd04911040;
                12'd3995: logsin <= 24'd04926010;
                12'd3996: logsin <= 24'd04941131;
                12'd3997: logsin <= 24'd04956404;
                12'd3998: logsin <= 24'd04971833;
                12'd3999: logsin <= 24'd04987422;
                12'd4000: logsin <= 24'd05003173;
                12'd4001: logsin <= 24'd05019090;
                12'd4002: logsin <= 24'd05035177;
                12'd4003: logsin <= 24'd05051436;
                12'd4004: logsin <= 24'd05067873;
                12'd4005: logsin <= 24'd05084490;
                12'd4006: logsin <= 24'd05101292;
                12'd4007: logsin <= 24'd05118283;
                12'd4008: logsin <= 24'd05135468;
                12'd4009: logsin <= 24'd05152850;
                12'd4010: logsin <= 24'd05170434;
                12'd4011: logsin <= 24'd05188225;
                12'd4012: logsin <= 24'd05206228;
                12'd4013: logsin <= 24'd05224448;
                12'd4014: logsin <= 24'd05242891;
                12'd4015: logsin <= 24'd05261562;
                12'd4016: logsin <= 24'd05280466;
                12'd4017: logsin <= 24'd05299609;
                12'd4018: logsin <= 24'd05318998;
                12'd4019: logsin <= 24'd05338639;
                12'd4020: logsin <= 24'd05358539;
                12'd4021: logsin <= 24'd05378704;
                12'd4022: logsin <= 24'd05399141;
                12'd4023: logsin <= 24'd05419859;
                12'd4024: logsin <= 24'd05440865;
                12'd4025: logsin <= 24'd05462167;
                12'd4026: logsin <= 24'd05483773;
                12'd4027: logsin <= 24'd05505693;
                12'd4028: logsin <= 24'd05527935;
                12'd4029: logsin <= 24'd05550509;
                12'd4030: logsin <= 24'd05573425;
                12'd4031: logsin <= 24'd05596694;
                12'd4032: logsin <= 24'd05620327;
                12'd4033: logsin <= 24'd05644335;
                12'd4034: logsin <= 24'd05668731;
                12'd4035: logsin <= 24'd05693527;
                12'd4036: logsin <= 24'd05718736;
                12'd4037: logsin <= 24'd05744372;
                12'd4038: logsin <= 24'd05770451;
                12'd4039: logsin <= 24'd05796987;
                12'd4040: logsin <= 24'd05823998;
                12'd4041: logsin <= 24'd05851499;
                12'd4042: logsin <= 24'd05879510;
                12'd4043: logsin <= 24'd05908050;
                12'd4044: logsin <= 24'd05937139;
                12'd4045: logsin <= 24'd05966799;
                12'd4046: logsin <= 24'd05997051;
                12'd4047: logsin <= 24'd06027922;
                12'd4048: logsin <= 24'd06059436;
                12'd4049: logsin <= 24'd06091620;
                12'd4050: logsin <= 24'd06124504;
                12'd4051: logsin <= 24'd06158120;
                12'd4052: logsin <= 24'd06192499;
                12'd4053: logsin <= 24'd06227678;
                12'd4054: logsin <= 24'd06263695;
                12'd4055: logsin <= 24'd06300591;
                12'd4056: logsin <= 24'd06338409;
                12'd4057: logsin <= 24'd06377198;
                12'd4058: logsin <= 24'd06417007;
                12'd4059: logsin <= 24'd06457893;
                12'd4060: logsin <= 24'd06499914;
                12'd4061: logsin <= 24'd06543137;
                12'd4062: logsin <= 24'd06587631;
                12'd4063: logsin <= 24'd06633474;
                12'd4064: logsin <= 24'd06680749;
                12'd4065: logsin <= 24'd06729550;
                12'd4066: logsin <= 24'd06779979;
                12'd4067: logsin <= 24'd06832146;
                12'd4068: logsin <= 24'd06886178;
                12'd4069: logsin <= 24'd06942211;
                12'd4070: logsin <= 24'd07000400;
                12'd4071: logsin <= 24'd07060917;
                12'd4072: logsin <= 24'd07123957;
                12'd4073: logsin <= 24'd07189738;
                12'd4074: logsin <= 24'd07258511;
                12'd4075: logsin <= 24'd07330560;
                12'd4076: logsin <= 24'd07406213;
                12'd4077: logsin <= 24'd07485850;
                12'd4078: logsin <= 24'd07569913;
                12'd4079: logsin <= 24'd07658924;
                12'd4080: logsin <= 24'd07753502;
                12'd4081: logsin <= 24'd07854390;
                12'd4082: logsin <= 24'd07962491;
                12'd4083: logsin <= 24'd08078914;
                12'd4084: logsin <= 24'd08205051;
                12'd4085: logsin <= 24'd08342670;
                12'd4086: logsin <= 24'd08494073;
                12'd4087: logsin <= 24'd08662332;
                12'd4088: logsin <= 24'd08851675;
                12'd4089: logsin <= 24'd09068154;
                12'd4090: logsin <= 24'd09320869;
                12'd4091: logsin <= 24'd09624438;
                12'd4092: logsin <= 24'd10004620;
                12'd4093: logsin <= 24'd10513627;
                12'd4094: logsin <= 24'd11286391;
                12'd4095: logsin <= 24'd12948345;
            endcase
        4'b01: //sine2xp 1/3 12/24-bit
            case (addr[15:4])
                12'd0000: logsin <= 24'd00000000;
                12'd0001: logsin <= 24'd00000000;
                12'd0002: logsin <= 24'd00000001;
                12'd0003: logsin <= 24'd00000002;
                12'd0004: logsin <= 24'd00000003;
                12'd0005: logsin <= 24'd00000005;
                12'd0006: logsin <= 24'd00000007;
                12'd0007: logsin <= 24'd00000009;
                12'd0008: logsin <= 24'd00000012;
                12'd0009: logsin <= 24'd00000015;
                12'd0010: logsin <= 24'd00000018;
                12'd0011: logsin <= 24'd00000022;
                12'd0012: logsin <= 24'd00000026;
                12'd0013: logsin <= 24'd00000030;
                12'd0014: logsin <= 24'd00000035;
                12'd0015: logsin <= 24'd00000040;
                12'd0016: logsin <= 24'd00000045;
                12'd0017: logsin <= 24'd00000051;
                12'd0018: logsin <= 24'd00000057;
                12'd0019: logsin <= 24'd00000063;
                12'd0020: logsin <= 24'd00000070;
                12'd0021: logsin <= 24'd00000077;
                12'd0022: logsin <= 24'd00000084;
                12'd0023: logsin <= 24'd00000092;
                12'd0024: logsin <= 24'd00000100;
                12'd0025: logsin <= 24'd00000108;
                12'd0026: logsin <= 24'd00000117;
                12'd0027: logsin <= 24'd00000126;
                12'd0028: logsin <= 24'd00000135;
                12'd0029: logsin <= 24'd00000145;
                12'd0030: logsin <= 24'd00000155;
                12'd0031: logsin <= 24'd00000165;
                12'd0032: logsin <= 24'd00000176;
                12'd0033: logsin <= 24'd00000187;
                12'd0034: logsin <= 24'd00000198;
                12'd0035: logsin <= 24'd00000210;
                12'd0036: logsin <= 24'd00000222;
                12'd0037: logsin <= 24'd00000234;
                12'd0038: logsin <= 24'd00000247;
                12'd0039: logsin <= 24'd00000260;
                12'd0040: logsin <= 24'd00000273;
                12'd0041: logsin <= 24'd00000287;
                12'd0042: logsin <= 24'd00000301;
                12'd0043: logsin <= 24'd00000315;
                12'd0044: logsin <= 24'd00000330;
                12'd0045: logsin <= 24'd00000345;
                12'd0046: logsin <= 24'd00000360;
                12'd0047: logsin <= 24'd00000376;
                12'd0048: logsin <= 24'd00000392;
                12'd0049: logsin <= 24'd00000408;
                12'd0050: logsin <= 24'd00000425;
                12'd0051: logsin <= 24'd00000442;
                12'd0052: logsin <= 24'd00000460;
                12'd0053: logsin <= 24'd00000477;
                12'd0054: logsin <= 24'd00000495;
                12'd0055: logsin <= 24'd00000514;
                12'd0056: logsin <= 24'd00000532;
                12'd0057: logsin <= 24'd00000551;
                12'd0058: logsin <= 24'd00000571;
                12'd0059: logsin <= 24'd00000590;
                12'd0060: logsin <= 24'd00000610;
                12'd0061: logsin <= 24'd00000631;
                12'd0062: logsin <= 24'd00000651;
                12'd0063: logsin <= 24'd00000672;
                12'd0064: logsin <= 24'd00000694;
                12'd0065: logsin <= 24'd00000716;
                12'd0066: logsin <= 24'd00000738;
                12'd0067: logsin <= 24'd00000760;
                12'd0068: logsin <= 24'd00000783;
                12'd0069: logsin <= 24'd00000806;
                12'd0070: logsin <= 24'd00000829;
                12'd0071: logsin <= 24'd00000853;
                12'd0072: logsin <= 24'd00000877;
                12'd0073: logsin <= 24'd00000901;
                12'd0074: logsin <= 24'd00000926;
                12'd0075: logsin <= 24'd00000951;
                12'd0076: logsin <= 24'd00000976;
                12'd0077: logsin <= 24'd00001002;
                12'd0078: logsin <= 24'd00001028;
                12'd0079: logsin <= 24'd00001054;
                12'd0080: logsin <= 24'd00001081;
                12'd0081: logsin <= 24'd00001108;
                12'd0082: logsin <= 24'd00001135;
                12'd0083: logsin <= 24'd00001163;
                12'd0084: logsin <= 24'd00001191;
                12'd0085: logsin <= 24'd00001219;
                12'd0086: logsin <= 24'd00001248;
                12'd0087: logsin <= 24'd00001277;
                12'd0088: logsin <= 24'd00001307;
                12'd0089: logsin <= 24'd00001336;
                12'd0090: logsin <= 24'd00001366;
                12'd0091: logsin <= 24'd00001397;
                12'd0092: logsin <= 24'd00001427;
                12'd0093: logsin <= 24'd00001458;
                12'd0094: logsin <= 24'd00001490;
                12'd0095: logsin <= 24'd00001522;
                12'd0096: logsin <= 24'd00001554;
                12'd0097: logsin <= 24'd00001586;
                12'd0098: logsin <= 24'd00001619;
                12'd0099: logsin <= 24'd00001652;
                12'd0100: logsin <= 24'd00001685;
                12'd0101: logsin <= 24'd00001719;
                12'd0102: logsin <= 24'd00001753;
                12'd0103: logsin <= 24'd00001787;
                12'd0104: logsin <= 24'd00001822;
                12'd0105: logsin <= 24'd00001857;
                12'd0106: logsin <= 24'd00001892;
                12'd0107: logsin <= 24'd00001928;
                12'd0108: logsin <= 24'd00001964;
                12'd0109: logsin <= 24'd00002000;
                12'd0110: logsin <= 24'd00002037;
                12'd0111: logsin <= 24'd00002074;
                12'd0112: logsin <= 24'd00002112;
                12'd0113: logsin <= 24'd00002149;
                12'd0114: logsin <= 24'd00002187;
                12'd0115: logsin <= 24'd00002226;
                12'd0116: logsin <= 24'd00002265;
                12'd0117: logsin <= 24'd00002304;
                12'd0118: logsin <= 24'd00002343;
                12'd0119: logsin <= 24'd00002383;
                12'd0120: logsin <= 24'd00002423;
                12'd0121: logsin <= 24'd00002463;
                12'd0122: logsin <= 24'd00002504;
                12'd0123: logsin <= 24'd00002545;
                12'd0124: logsin <= 24'd00002586;
                12'd0125: logsin <= 24'd00002628;
                12'd0126: logsin <= 24'd00002670;
                12'd0127: logsin <= 24'd00002712;
                12'd0128: logsin <= 24'd00002755;
                12'd0129: logsin <= 24'd00002798;
                12'd0130: logsin <= 24'd00002842;
                12'd0131: logsin <= 24'd00002885;
                12'd0132: logsin <= 24'd00002929;
                12'd0133: logsin <= 24'd00002974;
                12'd0134: logsin <= 24'd00003019;
                12'd0135: logsin <= 24'd00003064;
                12'd0136: logsin <= 24'd00003109;
                12'd0137: logsin <= 24'd00003155;
                12'd0138: logsin <= 24'd00003201;
                12'd0139: logsin <= 24'd00003247;
                12'd0140: logsin <= 24'd00003294;
                12'd0141: logsin <= 24'd00003341;
                12'd0142: logsin <= 24'd00003388;
                12'd0143: logsin <= 24'd00003436;
                12'd0144: logsin <= 24'd00003484;
                12'd0145: logsin <= 24'd00003533;
                12'd0146: logsin <= 24'd00003581;
                12'd0147: logsin <= 24'd00003630;
                12'd0148: logsin <= 24'd00003680;
                12'd0149: logsin <= 24'd00003730;
                12'd0150: logsin <= 24'd00003780;
                12'd0151: logsin <= 24'd00003830;
                12'd0152: logsin <= 24'd00003881;
                12'd0153: logsin <= 24'd00003932;
                12'd0154: logsin <= 24'd00003983;
                12'd0155: logsin <= 24'd00004035;
                12'd0156: logsin <= 24'd00004087;
                12'd0157: logsin <= 24'd00004139;
                12'd0158: logsin <= 24'd00004192;
                12'd0159: logsin <= 24'd00004245;
                12'd0160: logsin <= 24'd00004299;
                12'd0161: logsin <= 24'd00004352;
                12'd0162: logsin <= 24'd00004407;
                12'd0163: logsin <= 24'd00004461;
                12'd0164: logsin <= 24'd00004516;
                12'd0165: logsin <= 24'd00004571;
                12'd0166: logsin <= 24'd00004626;
                12'd0167: logsin <= 24'd00004682;
                12'd0168: logsin <= 24'd00004738;
                12'd0169: logsin <= 24'd00004794;
                12'd0170: logsin <= 24'd00004851;
                12'd0171: logsin <= 24'd00004908;
                12'd0172: logsin <= 24'd00004966;
                12'd0173: logsin <= 24'd00005023;
                12'd0174: logsin <= 24'd00005082;
                12'd0175: logsin <= 24'd00005140;
                12'd0176: logsin <= 24'd00005199;
                12'd0177: logsin <= 24'd00005258;
                12'd0178: logsin <= 24'd00005317;
                12'd0179: logsin <= 24'd00005377;
                12'd0180: logsin <= 24'd00005437;
                12'd0181: logsin <= 24'd00005498;
                12'd0182: logsin <= 24'd00005558;
                12'd0183: logsin <= 24'd00005619;
                12'd0184: logsin <= 24'd00005681;
                12'd0185: logsin <= 24'd00005743;
                12'd0186: logsin <= 24'd00005805;
                12'd0187: logsin <= 24'd00005867;
                12'd0188: logsin <= 24'd00005930;
                12'd0189: logsin <= 24'd00005993;
                12'd0190: logsin <= 24'd00006056;
                12'd0191: logsin <= 24'd00006120;
                12'd0192: logsin <= 24'd00006184;
                12'd0193: logsin <= 24'd00006249;
                12'd0194: logsin <= 24'd00006314;
                12'd0195: logsin <= 24'd00006379;
                12'd0196: logsin <= 24'd00006444;
                12'd0197: logsin <= 24'd00006510;
                12'd0198: logsin <= 24'd00006576;
                12'd0199: logsin <= 24'd00006642;
                12'd0200: logsin <= 24'd00006709;
                12'd0201: logsin <= 24'd00006776;
                12'd0202: logsin <= 24'd00006844;
                12'd0203: logsin <= 24'd00006911;
                12'd0204: logsin <= 24'd00006980;
                12'd0205: logsin <= 24'd00007048;
                12'd0206: logsin <= 24'd00007117;
                12'd0207: logsin <= 24'd00007186;
                12'd0208: logsin <= 24'd00007255;
                12'd0209: logsin <= 24'd00007325;
                12'd0210: logsin <= 24'd00007395;
                12'd0211: logsin <= 24'd00007466;
                12'd0212: logsin <= 24'd00007537;
                12'd0213: logsin <= 24'd00007608;
                12'd0214: logsin <= 24'd00007679;
                12'd0215: logsin <= 24'd00007751;
                12'd0216: logsin <= 24'd00007823;
                12'd0217: logsin <= 24'd00007896;
                12'd0218: logsin <= 24'd00007968;
                12'd0219: logsin <= 24'd00008041;
                12'd0220: logsin <= 24'd00008115;
                12'd0221: logsin <= 24'd00008189;
                12'd0222: logsin <= 24'd00008263;
                12'd0223: logsin <= 24'd00008337;
                12'd0224: logsin <= 24'd00008412;
                12'd0225: logsin <= 24'd00008487;
                12'd0226: logsin <= 24'd00008563;
                12'd0227: logsin <= 24'd00008638;
                12'd0228: logsin <= 24'd00008715;
                12'd0229: logsin <= 24'd00008791;
                12'd0230: logsin <= 24'd00008868;
                12'd0231: logsin <= 24'd00008945;
                12'd0232: logsin <= 24'd00009023;
                12'd0233: logsin <= 24'd00009100;
                12'd0234: logsin <= 24'd00009178;
                12'd0235: logsin <= 24'd00009257;
                12'd0236: logsin <= 24'd00009336;
                12'd0237: logsin <= 24'd00009415;
                12'd0238: logsin <= 24'd00009494;
                12'd0239: logsin <= 24'd00009574;
                12'd0240: logsin <= 24'd00009654;
                12'd0241: logsin <= 24'd00009735;
                12'd0242: logsin <= 24'd00009816;
                12'd0243: logsin <= 24'd00009897;
                12'd0244: logsin <= 24'd00009978;
                12'd0245: logsin <= 24'd00010060;
                12'd0246: logsin <= 24'd00010142;
                12'd0247: logsin <= 24'd00010225;
                12'd0248: logsin <= 24'd00010308;
                12'd0249: logsin <= 24'd00010391;
                12'd0250: logsin <= 24'd00010474;
                12'd0251: logsin <= 24'd00010558;
                12'd0252: logsin <= 24'd00010642;
                12'd0253: logsin <= 24'd00010727;
                12'd0254: logsin <= 24'd00010812;
                12'd0255: logsin <= 24'd00010897;
                12'd0256: logsin <= 24'd00010982;
                12'd0257: logsin <= 24'd00011068;
                12'd0258: logsin <= 24'd00011154;
                12'd0259: logsin <= 24'd00011241;
                12'd0260: logsin <= 24'd00011328;
                12'd0261: logsin <= 24'd00011415;
                12'd0262: logsin <= 24'd00011502;
                12'd0263: logsin <= 24'd00011590;
                12'd0264: logsin <= 24'd00011678;
                12'd0265: logsin <= 24'd00011767;
                12'd0266: logsin <= 24'd00011856;
                12'd0267: logsin <= 24'd00011945;
                12'd0268: logsin <= 24'd00012034;
                12'd0269: logsin <= 24'd00012124;
                12'd0270: logsin <= 24'd00012214;
                12'd0271: logsin <= 24'd00012305;
                12'd0272: logsin <= 24'd00012396;
                12'd0273: logsin <= 24'd00012487;
                12'd0274: logsin <= 24'd00012578;
                12'd0275: logsin <= 24'd00012670;
                12'd0276: logsin <= 24'd00012763;
                12'd0277: logsin <= 24'd00012855;
                12'd0278: logsin <= 24'd00012948;
                12'd0279: logsin <= 24'd00013041;
                12'd0280: logsin <= 24'd00013135;
                12'd0281: logsin <= 24'd00013228;
                12'd0282: logsin <= 24'd00013323;
                12'd0283: logsin <= 24'd00013417;
                12'd0284: logsin <= 24'd00013512;
                12'd0285: logsin <= 24'd00013607;
                12'd0286: logsin <= 24'd00013703;
                12'd0287: logsin <= 24'd00013799;
                12'd0288: logsin <= 24'd00013895;
                12'd0289: logsin <= 24'd00013991;
                12'd0290: logsin <= 24'd00014088;
                12'd0291: logsin <= 24'd00014186;
                12'd0292: logsin <= 24'd00014283;
                12'd0293: logsin <= 24'd00014381;
                12'd0294: logsin <= 24'd00014479;
                12'd0295: logsin <= 24'd00014578;
                12'd0296: logsin <= 24'd00014677;
                12'd0297: logsin <= 24'd00014776;
                12'd0298: logsin <= 24'd00014875;
                12'd0299: logsin <= 24'd00014975;
                12'd0300: logsin <= 24'd00015076;
                12'd0301: logsin <= 24'd00015176;
                12'd0302: logsin <= 24'd00015277;
                12'd0303: logsin <= 24'd00015378;
                12'd0304: logsin <= 24'd00015480;
                12'd0305: logsin <= 24'd00015582;
                12'd0306: logsin <= 24'd00015684;
                12'd0307: logsin <= 24'd00015787;
                12'd0308: logsin <= 24'd00015889;
                12'd0309: logsin <= 24'd00015993;
                12'd0310: logsin <= 24'd00016096;
                12'd0311: logsin <= 24'd00016200;
                12'd0312: logsin <= 24'd00016304;
                12'd0313: logsin <= 24'd00016409;
                12'd0314: logsin <= 24'd00016514;
                12'd0315: logsin <= 24'd00016619;
                12'd0316: logsin <= 24'd00016725;
                12'd0317: logsin <= 24'd00016831;
                12'd0318: logsin <= 24'd00016937;
                12'd0319: logsin <= 24'd00017043;
                12'd0320: logsin <= 24'd00017150;
                12'd0321: logsin <= 24'd00017258;
                12'd0322: logsin <= 24'd00017365;
                12'd0323: logsin <= 24'd00017473;
                12'd0324: logsin <= 24'd00017581;
                12'd0325: logsin <= 24'd00017690;
                12'd0326: logsin <= 24'd00017799;
                12'd0327: logsin <= 24'd00017908;
                12'd0328: logsin <= 24'd00018018;
                12'd0329: logsin <= 24'd00018128;
                12'd0330: logsin <= 24'd00018238;
                12'd0331: logsin <= 24'd00018349;
                12'd0332: logsin <= 24'd00018460;
                12'd0333: logsin <= 24'd00018571;
                12'd0334: logsin <= 24'd00018682;
                12'd0335: logsin <= 24'd00018794;
                12'd0336: logsin <= 24'd00018907;
                12'd0337: logsin <= 24'd00019019;
                12'd0338: logsin <= 24'd00019132;
                12'd0339: logsin <= 24'd00019246;
                12'd0340: logsin <= 24'd00019359;
                12'd0341: logsin <= 24'd00019473;
                12'd0342: logsin <= 24'd00019587;
                12'd0343: logsin <= 24'd00019702;
                12'd0344: logsin <= 24'd00019817;
                12'd0345: logsin <= 24'd00019932;
                12'd0346: logsin <= 24'd00020048;
                12'd0347: logsin <= 24'd00020164;
                12'd0348: logsin <= 24'd00020280;
                12'd0349: logsin <= 24'd00020397;
                12'd0350: logsin <= 24'd00020514;
                12'd0351: logsin <= 24'd00020631;
                12'd0352: logsin <= 24'd00020749;
                12'd0353: logsin <= 24'd00020867;
                12'd0354: logsin <= 24'd00020985;
                12'd0355: logsin <= 24'd00021104;
                12'd0356: logsin <= 24'd00021223;
                12'd0357: logsin <= 24'd00021342;
                12'd0358: logsin <= 24'd00021462;
                12'd0359: logsin <= 24'd00021582;
                12'd0360: logsin <= 24'd00021702;
                12'd0361: logsin <= 24'd00021823;
                12'd0362: logsin <= 24'd00021944;
                12'd0363: logsin <= 24'd00022065;
                12'd0364: logsin <= 24'd00022187;
                12'd0365: logsin <= 24'd00022309;
                12'd0366: logsin <= 24'd00022431;
                12'd0367: logsin <= 24'd00022554;
                12'd0368: logsin <= 24'd00022677;
                12'd0369: logsin <= 24'd00022800;
                12'd0370: logsin <= 24'd00022924;
                12'd0371: logsin <= 24'd00023048;
                12'd0372: logsin <= 24'd00023172;
                12'd0373: logsin <= 24'd00023297;
                12'd0374: logsin <= 24'd00023422;
                12'd0375: logsin <= 24'd00023547;
                12'd0376: logsin <= 24'd00023673;
                12'd0377: logsin <= 24'd00023799;
                12'd0378: logsin <= 24'd00023925;
                12'd0379: logsin <= 24'd00024052;
                12'd0380: logsin <= 24'd00024179;
                12'd0381: logsin <= 24'd00024306;
                12'd0382: logsin <= 24'd00024434;
                12'd0383: logsin <= 24'd00024562;
                12'd0384: logsin <= 24'd00024691;
                12'd0385: logsin <= 24'd00024819;
                12'd0386: logsin <= 24'd00024948;
                12'd0387: logsin <= 24'd00025078;
                12'd0388: logsin <= 24'd00025207;
                12'd0389: logsin <= 24'd00025338;
                12'd0390: logsin <= 24'd00025468;
                12'd0391: logsin <= 24'd00025599;
                12'd0392: logsin <= 24'd00025730;
                12'd0393: logsin <= 24'd00025861;
                12'd0394: logsin <= 24'd00025993;
                12'd0395: logsin <= 24'd00026125;
                12'd0396: logsin <= 24'd00026257;
                12'd0397: logsin <= 24'd00026390;
                12'd0398: logsin <= 24'd00026523;
                12'd0399: logsin <= 24'd00026657;
                12'd0400: logsin <= 24'd00026790;
                12'd0401: logsin <= 24'd00026924;
                12'd0402: logsin <= 24'd00027059;
                12'd0403: logsin <= 24'd00027194;
                12'd0404: logsin <= 24'd00027329;
                12'd0405: logsin <= 24'd00027464;
                12'd0406: logsin <= 24'd00027600;
                12'd0407: logsin <= 24'd00027736;
                12'd0408: logsin <= 24'd00027872;
                12'd0409: logsin <= 24'd00028009;
                12'd0410: logsin <= 24'd00028146;
                12'd0411: logsin <= 24'd00028284;
                12'd0412: logsin <= 24'd00028421;
                12'd0413: logsin <= 24'd00028560;
                12'd0414: logsin <= 24'd00028698;
                12'd0415: logsin <= 24'd00028837;
                12'd0416: logsin <= 24'd00028976;
                12'd0417: logsin <= 24'd00029115;
                12'd0418: logsin <= 24'd00029255;
                12'd0419: logsin <= 24'd00029395;
                12'd0420: logsin <= 24'd00029536;
                12'd0421: logsin <= 24'd00029676;
                12'd0422: logsin <= 24'd00029818;
                12'd0423: logsin <= 24'd00029959;
                12'd0424: logsin <= 24'd00030101;
                12'd0425: logsin <= 24'd00030243;
                12'd0426: logsin <= 24'd00030386;
                12'd0427: logsin <= 24'd00030528;
                12'd0428: logsin <= 24'd00030671;
                12'd0429: logsin <= 24'd00030815;
                12'd0430: logsin <= 24'd00030959;
                12'd0431: logsin <= 24'd00031103;
                12'd0432: logsin <= 24'd00031247;
                12'd0433: logsin <= 24'd00031392;
                12'd0434: logsin <= 24'd00031537;
                12'd0435: logsin <= 24'd00031683;
                12'd0436: logsin <= 24'd00031829;
                12'd0437: logsin <= 24'd00031975;
                12'd0438: logsin <= 24'd00032121;
                12'd0439: logsin <= 24'd00032268;
                12'd0440: logsin <= 24'd00032415;
                12'd0441: logsin <= 24'd00032563;
                12'd0442: logsin <= 24'd00032711;
                12'd0443: logsin <= 24'd00032859;
                12'd0444: logsin <= 24'd00033008;
                12'd0445: logsin <= 24'd00033156;
                12'd0446: logsin <= 24'd00033306;
                12'd0447: logsin <= 24'd00033455;
                12'd0448: logsin <= 24'd00033605;
                12'd0449: logsin <= 24'd00033755;
                12'd0450: logsin <= 24'd00033906;
                12'd0451: logsin <= 24'd00034057;
                12'd0452: logsin <= 24'd00034208;
                12'd0453: logsin <= 24'd00034359;
                12'd0454: logsin <= 24'd00034511;
                12'd0455: logsin <= 24'd00034663;
                12'd0456: logsin <= 24'd00034816;
                12'd0457: logsin <= 24'd00034969;
                12'd0458: logsin <= 24'd00035122;
                12'd0459: logsin <= 24'd00035276;
                12'd0460: logsin <= 24'd00035430;
                12'd0461: logsin <= 24'd00035584;
                12'd0462: logsin <= 24'd00035738;
                12'd0463: logsin <= 24'd00035893;
                12'd0464: logsin <= 24'd00036049;
                12'd0465: logsin <= 24'd00036204;
                12'd0466: logsin <= 24'd00036360;
                12'd0467: logsin <= 24'd00036516;
                12'd0468: logsin <= 24'd00036673;
                12'd0469: logsin <= 24'd00036830;
                12'd0470: logsin <= 24'd00036987;
                12'd0471: logsin <= 24'd00037145;
                12'd0472: logsin <= 24'd00037303;
                12'd0473: logsin <= 24'd00037461;
                12'd0474: logsin <= 24'd00037620;
                12'd0475: logsin <= 24'd00037779;
                12'd0476: logsin <= 24'd00037938;
                12'd0477: logsin <= 24'd00038097;
                12'd0478: logsin <= 24'd00038257;
                12'd0479: logsin <= 24'd00038418;
                12'd0480: logsin <= 24'd00038578;
                12'd0481: logsin <= 24'd00038739;
                12'd0482: logsin <= 24'd00038901;
                12'd0483: logsin <= 24'd00039062;
                12'd0484: logsin <= 24'd00039224;
                12'd0485: logsin <= 24'd00039386;
                12'd0486: logsin <= 24'd00039549;
                12'd0487: logsin <= 24'd00039712;
                12'd0488: logsin <= 24'd00039875;
                12'd0489: logsin <= 24'd00040039;
                12'd0490: logsin <= 24'd00040203;
                12'd0491: logsin <= 24'd00040367;
                12'd0492: logsin <= 24'd00040532;
                12'd0493: logsin <= 24'd00040697;
                12'd0494: logsin <= 24'd00040862;
                12'd0495: logsin <= 24'd00041028;
                12'd0496: logsin <= 24'd00041194;
                12'd0497: logsin <= 24'd00041360;
                12'd0498: logsin <= 24'd00041527;
                12'd0499: logsin <= 24'd00041694;
                12'd0500: logsin <= 24'd00041862;
                12'd0501: logsin <= 24'd00042029;
                12'd0502: logsin <= 24'd00042197;
                12'd0503: logsin <= 24'd00042366;
                12'd0504: logsin <= 24'd00042534;
                12'd0505: logsin <= 24'd00042703;
                12'd0506: logsin <= 24'd00042873;
                12'd0507: logsin <= 24'd00043042;
                12'd0508: logsin <= 24'd00043213;
                12'd0509: logsin <= 24'd00043383;
                12'd0510: logsin <= 24'd00043554;
                12'd0511: logsin <= 24'd00043725;
                12'd0512: logsin <= 24'd00043896;
                12'd0513: logsin <= 24'd00044068;
                12'd0514: logsin <= 24'd00044240;
                12'd0515: logsin <= 24'd00044412;
                12'd0516: logsin <= 24'd00044585;
                12'd0517: logsin <= 24'd00044758;
                12'd0518: logsin <= 24'd00044932;
                12'd0519: logsin <= 24'd00045105;
                12'd0520: logsin <= 24'd00045279;
                12'd0521: logsin <= 24'd00045454;
                12'd0522: logsin <= 24'd00045629;
                12'd0523: logsin <= 24'd00045804;
                12'd0524: logsin <= 24'd00045979;
                12'd0525: logsin <= 24'd00046155;
                12'd0526: logsin <= 24'd00046331;
                12'd0527: logsin <= 24'd00046508;
                12'd0528: logsin <= 24'd00046684;
                12'd0529: logsin <= 24'd00046861;
                12'd0530: logsin <= 24'd00047039;
                12'd0531: logsin <= 24'd00047217;
                12'd0532: logsin <= 24'd00047395;
                12'd0533: logsin <= 24'd00047573;
                12'd0534: logsin <= 24'd00047752;
                12'd0535: logsin <= 24'd00047931;
                12'd0536: logsin <= 24'd00048111;
                12'd0537: logsin <= 24'd00048291;
                12'd0538: logsin <= 24'd00048471;
                12'd0539: logsin <= 24'd00048651;
                12'd0540: logsin <= 24'd00048832;
                12'd0541: logsin <= 24'd00049013;
                12'd0542: logsin <= 24'd00049195;
                12'd0543: logsin <= 24'd00049377;
                12'd0544: logsin <= 24'd00049559;
                12'd0545: logsin <= 24'd00049741;
                12'd0546: logsin <= 24'd00049924;
                12'd0547: logsin <= 24'd00050107;
                12'd0548: logsin <= 24'd00050291;
                12'd0549: logsin <= 24'd00050475;
                12'd0550: logsin <= 24'd00050659;
                12'd0551: logsin <= 24'd00050844;
                12'd0552: logsin <= 24'd00051028;
                12'd0553: logsin <= 24'd00051214;
                12'd0554: logsin <= 24'd00051399;
                12'd0555: logsin <= 24'd00051585;
                12'd0556: logsin <= 24'd00051771;
                12'd0557: logsin <= 24'd00051958;
                12'd0558: logsin <= 24'd00052145;
                12'd0559: logsin <= 24'd00052332;
                12'd0560: logsin <= 24'd00052520;
                12'd0561: logsin <= 24'd00052708;
                12'd0562: logsin <= 24'd00052896;
                12'd0563: logsin <= 24'd00053084;
                12'd0564: logsin <= 24'd00053273;
                12'd0565: logsin <= 24'd00053463;
                12'd0566: logsin <= 24'd00053652;
                12'd0567: logsin <= 24'd00053842;
                12'd0568: logsin <= 24'd00054032;
                12'd0569: logsin <= 24'd00054223;
                12'd0570: logsin <= 24'd00054414;
                12'd0571: logsin <= 24'd00054605;
                12'd0572: logsin <= 24'd00054797;
                12'd0573: logsin <= 24'd00054989;
                12'd0574: logsin <= 24'd00055181;
                12'd0575: logsin <= 24'd00055374;
                12'd0576: logsin <= 24'd00055567;
                12'd0577: logsin <= 24'd00055760;
                12'd0578: logsin <= 24'd00055954;
                12'd0579: logsin <= 24'd00056148;
                12'd0580: logsin <= 24'd00056342;
                12'd0581: logsin <= 24'd00056537;
                12'd0582: logsin <= 24'd00056732;
                12'd0583: logsin <= 24'd00056927;
                12'd0584: logsin <= 24'd00057123;
                12'd0585: logsin <= 24'd00057319;
                12'd0586: logsin <= 24'd00057515;
                12'd0587: logsin <= 24'd00057712;
                12'd0588: logsin <= 24'd00057909;
                12'd0589: logsin <= 24'd00058106;
                12'd0590: logsin <= 24'd00058304;
                12'd0591: logsin <= 24'd00058502;
                12'd0592: logsin <= 24'd00058700;
                12'd0593: logsin <= 24'd00058899;
                12'd0594: logsin <= 24'd00059098;
                12'd0595: logsin <= 24'd00059298;
                12'd0596: logsin <= 24'd00059497;
                12'd0597: logsin <= 24'd00059697;
                12'd0598: logsin <= 24'd00059898;
                12'd0599: logsin <= 24'd00060099;
                12'd0600: logsin <= 24'd00060300;
                12'd0601: logsin <= 24'd00060501;
                12'd0602: logsin <= 24'd00060703;
                12'd0603: logsin <= 24'd00060905;
                12'd0604: logsin <= 24'd00061107;
                12'd0605: logsin <= 24'd00061310;
                12'd0606: logsin <= 24'd00061513;
                12'd0607: logsin <= 24'd00061717;
                12'd0608: logsin <= 24'd00061921;
                12'd0609: logsin <= 24'd00062125;
                12'd0610: logsin <= 24'd00062329;
                12'd0611: logsin <= 24'd00062534;
                12'd0612: logsin <= 24'd00062739;
                12'd0613: logsin <= 24'd00062945;
                12'd0614: logsin <= 24'd00063150;
                12'd0615: logsin <= 24'd00063357;
                12'd0616: logsin <= 24'd00063563;
                12'd0617: logsin <= 24'd00063770;
                12'd0618: logsin <= 24'd00063977;
                12'd0619: logsin <= 24'd00064185;
                12'd0620: logsin <= 24'd00064392;
                12'd0621: logsin <= 24'd00064601;
                12'd0622: logsin <= 24'd00064809;
                12'd0623: logsin <= 24'd00065018;
                12'd0624: logsin <= 24'd00065227;
                12'd0625: logsin <= 24'd00065437;
                12'd0626: logsin <= 24'd00065647;
                12'd0627: logsin <= 24'd00065857;
                12'd0628: logsin <= 24'd00066067;
                12'd0629: logsin <= 24'd00066278;
                12'd0630: logsin <= 24'd00066489;
                12'd0631: logsin <= 24'd00066701;
                12'd0632: logsin <= 24'd00066913;
                12'd0633: logsin <= 24'd00067125;
                12'd0634: logsin <= 24'd00067338;
                12'd0635: logsin <= 24'd00067551;
                12'd0636: logsin <= 24'd00067764;
                12'd0637: logsin <= 24'd00067977;
                12'd0638: logsin <= 24'd00068191;
                12'd0639: logsin <= 24'd00068406;
                12'd0640: logsin <= 24'd00068620;
                12'd0641: logsin <= 24'd00068835;
                12'd0642: logsin <= 24'd00069051;
                12'd0643: logsin <= 24'd00069266;
                12'd0644: logsin <= 24'd00069482;
                12'd0645: logsin <= 24'd00069698;
                12'd0646: logsin <= 24'd00069915;
                12'd0647: logsin <= 24'd00070132;
                12'd0648: logsin <= 24'd00070349;
                12'd0649: logsin <= 24'd00070567;
                12'd0650: logsin <= 24'd00070785;
                12'd0651: logsin <= 24'd00071003;
                12'd0652: logsin <= 24'd00071222;
                12'd0653: logsin <= 24'd00071441;
                12'd0654: logsin <= 24'd00071660;
                12'd0655: logsin <= 24'd00071880;
                12'd0656: logsin <= 24'd00072100;
                12'd0657: logsin <= 24'd00072320;
                12'd0658: logsin <= 24'd00072541;
                12'd0659: logsin <= 24'd00072762;
                12'd0660: logsin <= 24'd00072984;
                12'd0661: logsin <= 24'd00073205;
                12'd0662: logsin <= 24'd00073427;
                12'd0663: logsin <= 24'd00073650;
                12'd0664: logsin <= 24'd00073872;
                12'd0665: logsin <= 24'd00074096;
                12'd0666: logsin <= 24'd00074319;
                12'd0667: logsin <= 24'd00074543;
                12'd0668: logsin <= 24'd00074767;
                12'd0669: logsin <= 24'd00074991;
                12'd0670: logsin <= 24'd00075216;
                12'd0671: logsin <= 24'd00075441;
                12'd0672: logsin <= 24'd00075667;
                12'd0673: logsin <= 24'd00075892;
                12'd0674: logsin <= 24'd00076118;
                12'd0675: logsin <= 24'd00076345;
                12'd0676: logsin <= 24'd00076572;
                12'd0677: logsin <= 24'd00076799;
                12'd0678: logsin <= 24'd00077026;
                12'd0679: logsin <= 24'd00077254;
                12'd0680: logsin <= 24'd00077482;
                12'd0681: logsin <= 24'd00077711;
                12'd0682: logsin <= 24'd00077940;
                12'd0683: logsin <= 24'd00078169;
                12'd0684: logsin <= 24'd00078398;
                12'd0685: logsin <= 24'd00078628;
                12'd0686: logsin <= 24'd00078858;
                12'd0687: logsin <= 24'd00079089;
                12'd0688: logsin <= 24'd00079320;
                12'd0689: logsin <= 24'd00079551;
                12'd0690: logsin <= 24'd00079783;
                12'd0691: logsin <= 24'd00080014;
                12'd0692: logsin <= 24'd00080247;
                12'd0693: logsin <= 24'd00080479;
                12'd0694: logsin <= 24'd00080712;
                12'd0695: logsin <= 24'd00080945;
                12'd0696: logsin <= 24'd00081179;
                12'd0697: logsin <= 24'd00081413;
                12'd0698: logsin <= 24'd00081647;
                12'd0699: logsin <= 24'd00081882;
                12'd0700: logsin <= 24'd00082117;
                12'd0701: logsin <= 24'd00082352;
                12'd0702: logsin <= 24'd00082588;
                12'd0703: logsin <= 24'd00082824;
                12'd0704: logsin <= 24'd00083060;
                12'd0705: logsin <= 24'd00083296;
                12'd0706: logsin <= 24'd00083533;
                12'd0707: logsin <= 24'd00083771;
                12'd0708: logsin <= 24'd00084008;
                12'd0709: logsin <= 24'd00084246;
                12'd0710: logsin <= 24'd00084485;
                12'd0711: logsin <= 24'd00084723;
                12'd0712: logsin <= 24'd00084962;
                12'd0713: logsin <= 24'd00085202;
                12'd0714: logsin <= 24'd00085441;
                12'd0715: logsin <= 24'd00085682;
                12'd0716: logsin <= 24'd00085922;
                12'd0717: logsin <= 24'd00086163;
                12'd0718: logsin <= 24'd00086404;
                12'd0719: logsin <= 24'd00086645;
                12'd0720: logsin <= 24'd00086887;
                12'd0721: logsin <= 24'd00087129;
                12'd0722: logsin <= 24'd00087371;
                12'd0723: logsin <= 24'd00087614;
                12'd0724: logsin <= 24'd00087857;
                12'd0725: logsin <= 24'd00088100;
                12'd0726: logsin <= 24'd00088344;
                12'd0727: logsin <= 24'd00088588;
                12'd0728: logsin <= 24'd00088833;
                12'd0729: logsin <= 24'd00089078;
                12'd0730: logsin <= 24'd00089323;
                12'd0731: logsin <= 24'd00089568;
                12'd0732: logsin <= 24'd00089814;
                12'd0733: logsin <= 24'd00090060;
                12'd0734: logsin <= 24'd00090307;
                12'd0735: logsin <= 24'd00090553;
                12'd0736: logsin <= 24'd00090801;
                12'd0737: logsin <= 24'd00091048;
                12'd0738: logsin <= 24'd00091296;
                12'd0739: logsin <= 24'd00091544;
                12'd0740: logsin <= 24'd00091793;
                12'd0741: logsin <= 24'd00092041;
                12'd0742: logsin <= 24'd00092291;
                12'd0743: logsin <= 24'd00092540;
                12'd0744: logsin <= 24'd00092790;
                12'd0745: logsin <= 24'd00093040;
                12'd0746: logsin <= 24'd00093291;
                12'd0747: logsin <= 24'd00093542;
                12'd0748: logsin <= 24'd00093793;
                12'd0749: logsin <= 24'd00094045;
                12'd0750: logsin <= 24'd00094296;
                12'd0751: logsin <= 24'd00094549;
                12'd0752: logsin <= 24'd00094801;
                12'd0753: logsin <= 24'd00095054;
                12'd0754: logsin <= 24'd00095308;
                12'd0755: logsin <= 24'd00095561;
                12'd0756: logsin <= 24'd00095815;
                12'd0757: logsin <= 24'd00096069;
                12'd0758: logsin <= 24'd00096324;
                12'd0759: logsin <= 24'd00096579;
                12'd0760: logsin <= 24'd00096834;
                12'd0761: logsin <= 24'd00097090;
                12'd0762: logsin <= 24'd00097346;
                12'd0763: logsin <= 24'd00097602;
                12'd0764: logsin <= 24'd00097859;
                12'd0765: logsin <= 24'd00098116;
                12'd0766: logsin <= 24'd00098373;
                12'd0767: logsin <= 24'd00098631;
                12'd0768: logsin <= 24'd00098889;
                12'd0769: logsin <= 24'd00099148;
                12'd0770: logsin <= 24'd00099406;
                12'd0771: logsin <= 24'd00099665;
                12'd0772: logsin <= 24'd00099925;
                12'd0773: logsin <= 24'd00100184;
                12'd0774: logsin <= 24'd00100445;
                12'd0775: logsin <= 24'd00100705;
                12'd0776: logsin <= 24'd00100966;
                12'd0777: logsin <= 24'd00101227;
                12'd0778: logsin <= 24'd00101488;
                12'd0779: logsin <= 24'd00101750;
                12'd0780: logsin <= 24'd00102012;
                12'd0781: logsin <= 24'd00102275;
                12'd0782: logsin <= 24'd00102537;
                12'd0783: logsin <= 24'd00102801;
                12'd0784: logsin <= 24'd00103064;
                12'd0785: logsin <= 24'd00103328;
                12'd0786: logsin <= 24'd00103592;
                12'd0787: logsin <= 24'd00103857;
                12'd0788: logsin <= 24'd00104121;
                12'd0789: logsin <= 24'd00104387;
                12'd0790: logsin <= 24'd00104652;
                12'd0791: logsin <= 24'd00104918;
                12'd0792: logsin <= 24'd00105184;
                12'd0793: logsin <= 24'd00105451;
                12'd0794: logsin <= 24'd00105718;
                12'd0795: logsin <= 24'd00105985;
                12'd0796: logsin <= 24'd00106252;
                12'd0797: logsin <= 24'd00106520;
                12'd0798: logsin <= 24'd00106789;
                12'd0799: logsin <= 24'd00107057;
                12'd0800: logsin <= 24'd00107326;
                12'd0801: logsin <= 24'd00107595;
                12'd0802: logsin <= 24'd00107865;
                12'd0803: logsin <= 24'd00108135;
                12'd0804: logsin <= 24'd00108405;
                12'd0805: logsin <= 24'd00108676;
                12'd0806: logsin <= 24'd00108947;
                12'd0807: logsin <= 24'd00109218;
                12'd0808: logsin <= 24'd00109490;
                12'd0809: logsin <= 24'd00109762;
                12'd0810: logsin <= 24'd00110034;
                12'd0811: logsin <= 24'd00110307;
                12'd0812: logsin <= 24'd00110580;
                12'd0813: logsin <= 24'd00110853;
                12'd0814: logsin <= 24'd00111127;
                12'd0815: logsin <= 24'd00111401;
                12'd0816: logsin <= 24'd00111675;
                12'd0817: logsin <= 24'd00111950;
                12'd0818: logsin <= 24'd00112225;
                12'd0819: logsin <= 24'd00112501;
                12'd0820: logsin <= 24'd00112776;
                12'd0821: logsin <= 24'd00113053;
                12'd0822: logsin <= 24'd00113329;
                12'd0823: logsin <= 24'd00113606;
                12'd0824: logsin <= 24'd00113883;
                12'd0825: logsin <= 24'd00114160;
                12'd0826: logsin <= 24'd00114438;
                12'd0827: logsin <= 24'd00114716;
                12'd0828: logsin <= 24'd00114995;
                12'd0829: logsin <= 24'd00115274;
                12'd0830: logsin <= 24'd00115553;
                12'd0831: logsin <= 24'd00115832;
                12'd0832: logsin <= 24'd00116112;
                12'd0833: logsin <= 24'd00116392;
                12'd0834: logsin <= 24'd00116673;
                12'd0835: logsin <= 24'd00116954;
                12'd0836: logsin <= 24'd00117235;
                12'd0837: logsin <= 24'd00117516;
                12'd0838: logsin <= 24'd00117798;
                12'd0839: logsin <= 24'd00118081;
                12'd0840: logsin <= 24'd00118363;
                12'd0841: logsin <= 24'd00118646;
                12'd0842: logsin <= 24'd00118929;
                12'd0843: logsin <= 24'd00119213;
                12'd0844: logsin <= 24'd00119497;
                12'd0845: logsin <= 24'd00119781;
                12'd0846: logsin <= 24'd00120066;
                12'd0847: logsin <= 24'd00120351;
                12'd0848: logsin <= 24'd00120636;
                12'd0849: logsin <= 24'd00120922;
                12'd0850: logsin <= 24'd00121208;
                12'd0851: logsin <= 24'd00121494;
                12'd0852: logsin <= 24'd00121781;
                12'd0853: logsin <= 24'd00122068;
                12'd0854: logsin <= 24'd00122355;
                12'd0855: logsin <= 24'd00122643;
                12'd0856: logsin <= 24'd00122931;
                12'd0857: logsin <= 24'd00123219;
                12'd0858: logsin <= 24'd00123508;
                12'd0859: logsin <= 24'd00123797;
                12'd0860: logsin <= 24'd00124086;
                12'd0861: logsin <= 24'd00124376;
                12'd0862: logsin <= 24'd00124666;
                12'd0863: logsin <= 24'd00124957;
                12'd0864: logsin <= 24'd00125247;
                12'd0865: logsin <= 24'd00125538;
                12'd0866: logsin <= 24'd00125830;
                12'd0867: logsin <= 24'd00126122;
                12'd0868: logsin <= 24'd00126414;
                12'd0869: logsin <= 24'd00126706;
                12'd0870: logsin <= 24'd00126999;
                12'd0871: logsin <= 24'd00127292;
                12'd0872: logsin <= 24'd00127586;
                12'd0873: logsin <= 24'd00127880;
                12'd0874: logsin <= 24'd00128174;
                12'd0875: logsin <= 24'd00128468;
                12'd0876: logsin <= 24'd00128763;
                12'd0877: logsin <= 24'd00129058;
                12'd0878: logsin <= 24'd00129354;
                12'd0879: logsin <= 24'd00129650;
                12'd0880: logsin <= 24'd00129946;
                12'd0881: logsin <= 24'd00130243;
                12'd0882: logsin <= 24'd00130540;
                12'd0883: logsin <= 24'd00130837;
                12'd0884: logsin <= 24'd00131134;
                12'd0885: logsin <= 24'd00131432;
                12'd0886: logsin <= 24'd00131731;
                12'd0887: logsin <= 24'd00132029;
                12'd0888: logsin <= 24'd00132328;
                12'd0889: logsin <= 24'd00132628;
                12'd0890: logsin <= 24'd00132927;
                12'd0891: logsin <= 24'd00133227;
                12'd0892: logsin <= 24'd00133528;
                12'd0893: logsin <= 24'd00133828;
                12'd0894: logsin <= 24'd00134129;
                12'd0895: logsin <= 24'd00134431;
                12'd0896: logsin <= 24'd00134732;
                12'd0897: logsin <= 24'd00135034;
                12'd0898: logsin <= 24'd00135337;
                12'd0899: logsin <= 24'd00135640;
                12'd0900: logsin <= 24'd00135943;
                12'd0901: logsin <= 24'd00136246;
                12'd0902: logsin <= 24'd00136550;
                12'd0903: logsin <= 24'd00136854;
                12'd0904: logsin <= 24'd00137158;
                12'd0905: logsin <= 24'd00137463;
                12'd0906: logsin <= 24'd00137768;
                12'd0907: logsin <= 24'd00138074;
                12'd0908: logsin <= 24'd00138380;
                12'd0909: logsin <= 24'd00138686;
                12'd0910: logsin <= 24'd00138992;
                12'd0911: logsin <= 24'd00139299;
                12'd0912: logsin <= 24'd00139606;
                12'd0913: logsin <= 24'd00139914;
                12'd0914: logsin <= 24'd00140222;
                12'd0915: logsin <= 24'd00140530;
                12'd0916: logsin <= 24'd00140838;
                12'd0917: logsin <= 24'd00141147;
                12'd0918: logsin <= 24'd00141457;
                12'd0919: logsin <= 24'd00141766;
                12'd0920: logsin <= 24'd00142076;
                12'd0921: logsin <= 24'd00142386;
                12'd0922: logsin <= 24'd00142697;
                12'd0923: logsin <= 24'd00143008;
                12'd0924: logsin <= 24'd00143319;
                12'd0925: logsin <= 24'd00143631;
                12'd0926: logsin <= 24'd00143943;
                12'd0927: logsin <= 24'd00144255;
                12'd0928: logsin <= 24'd00144568;
                12'd0929: logsin <= 24'd00144881;
                12'd0930: logsin <= 24'd00145194;
                12'd0931: logsin <= 24'd00145508;
                12'd0932: logsin <= 24'd00145822;
                12'd0933: logsin <= 24'd00146136;
                12'd0934: logsin <= 24'd00146451;
                12'd0935: logsin <= 24'd00146766;
                12'd0936: logsin <= 24'd00147082;
                12'd0937: logsin <= 24'd00147397;
                12'd0938: logsin <= 24'd00147713;
                12'd0939: logsin <= 24'd00148030;
                12'd0940: logsin <= 24'd00148347;
                12'd0941: logsin <= 24'd00148664;
                12'd0942: logsin <= 24'd00148981;
                12'd0943: logsin <= 24'd00149299;
                12'd0944: logsin <= 24'd00149617;
                12'd0945: logsin <= 24'd00149936;
                12'd0946: logsin <= 24'd00150255;
                12'd0947: logsin <= 24'd00150574;
                12'd0948: logsin <= 24'd00150893;
                12'd0949: logsin <= 24'd00151213;
                12'd0950: logsin <= 24'd00151533;
                12'd0951: logsin <= 24'd00151854;
                12'd0952: logsin <= 24'd00152175;
                12'd0953: logsin <= 24'd00152496;
                12'd0954: logsin <= 24'd00152818;
                12'd0955: logsin <= 24'd00153139;
                12'd0956: logsin <= 24'd00153462;
                12'd0957: logsin <= 24'd00153784;
                12'd0958: logsin <= 24'd00154107;
                12'd0959: logsin <= 24'd00154431;
                12'd0960: logsin <= 24'd00154754;
                12'd0961: logsin <= 24'd00155078;
                12'd0962: logsin <= 24'd00155403;
                12'd0963: logsin <= 24'd00155727;
                12'd0964: logsin <= 24'd00156052;
                12'd0965: logsin <= 24'd00156378;
                12'd0966: logsin <= 24'd00156703;
                12'd0967: logsin <= 24'd00157029;
                12'd0968: logsin <= 24'd00157356;
                12'd0969: logsin <= 24'd00157682;
                12'd0970: logsin <= 24'd00158009;
                12'd0971: logsin <= 24'd00158337;
                12'd0972: logsin <= 24'd00158665;
                12'd0973: logsin <= 24'd00158993;
                12'd0974: logsin <= 24'd00159321;
                12'd0975: logsin <= 24'd00159650;
                12'd0976: logsin <= 24'd00159979;
                12'd0977: logsin <= 24'd00160309;
                12'd0978: logsin <= 24'd00160638;
                12'd0979: logsin <= 24'd00160969;
                12'd0980: logsin <= 24'd00161299;
                12'd0981: logsin <= 24'd00161630;
                12'd0982: logsin <= 24'd00161961;
                12'd0983: logsin <= 24'd00162293;
                12'd0984: logsin <= 24'd00162625;
                12'd0985: logsin <= 24'd00162957;
                12'd0986: logsin <= 24'd00163289;
                12'd0987: logsin <= 24'd00163622;
                12'd0988: logsin <= 24'd00163955;
                12'd0989: logsin <= 24'd00164289;
                12'd0990: logsin <= 24'd00164623;
                12'd0991: logsin <= 24'd00164957;
                12'd0992: logsin <= 24'd00165292;
                12'd0993: logsin <= 24'd00165627;
                12'd0994: logsin <= 24'd00165962;
                12'd0995: logsin <= 24'd00166298;
                12'd0996: logsin <= 24'd00166634;
                12'd0997: logsin <= 24'd00166970;
                12'd0998: logsin <= 24'd00167307;
                12'd0999: logsin <= 24'd00167644;
                12'd1000: logsin <= 24'd00167981;
                12'd1001: logsin <= 24'd00168319;
                12'd1002: logsin <= 24'd00168657;
                12'd1003: logsin <= 24'd00168996;
                12'd1004: logsin <= 24'd00169334;
                12'd1005: logsin <= 24'd00169673;
                12'd1006: logsin <= 24'd00170013;
                12'd1007: logsin <= 24'd00170353;
                12'd1008: logsin <= 24'd00170693;
                12'd1009: logsin <= 24'd00171033;
                12'd1010: logsin <= 24'd00171374;
                12'd1011: logsin <= 24'd00171715;
                12'd1012: logsin <= 24'd00172057;
                12'd1013: logsin <= 24'd00172398;
                12'd1014: logsin <= 24'd00172741;
                12'd1015: logsin <= 24'd00173083;
                12'd1016: logsin <= 24'd00173426;
                12'd1017: logsin <= 24'd00173769;
                12'd1018: logsin <= 24'd00174113;
                12'd1019: logsin <= 24'd00174457;
                12'd1020: logsin <= 24'd00174801;
                12'd1021: logsin <= 24'd00175146;
                12'd1022: logsin <= 24'd00175491;
                12'd1023: logsin <= 24'd00175836;
                12'd1024: logsin <= 24'd00176181;
                12'd1025: logsin <= 24'd00176527;
                12'd1026: logsin <= 24'd00176874;
                12'd1027: logsin <= 24'd00177220;
                12'd1028: logsin <= 24'd00177567;
                12'd1029: logsin <= 24'd00177915;
                12'd1030: logsin <= 24'd00178262;
                12'd1031: logsin <= 24'd00178611;
                12'd1032: logsin <= 24'd00178959;
                12'd1033: logsin <= 24'd00179308;
                12'd1034: logsin <= 24'd00179657;
                12'd1035: logsin <= 24'd00180006;
                12'd1036: logsin <= 24'd00180356;
                12'd1037: logsin <= 24'd00180706;
                12'd1038: logsin <= 24'd00181056;
                12'd1039: logsin <= 24'd00181407;
                12'd1040: logsin <= 24'd00181758;
                12'd1041: logsin <= 24'd00182110;
                12'd1042: logsin <= 24'd00182462;
                12'd1043: logsin <= 24'd00182814;
                12'd1044: logsin <= 24'd00183166;
                12'd1045: logsin <= 24'd00183519;
                12'd1046: logsin <= 24'd00183872;
                12'd1047: logsin <= 24'd00184226;
                12'd1048: logsin <= 24'd00184580;
                12'd1049: logsin <= 24'd00184934;
                12'd1050: logsin <= 24'd00185289;
                12'd1051: logsin <= 24'd00185644;
                12'd1052: logsin <= 24'd00185999;
                12'd1053: logsin <= 24'd00186354;
                12'd1054: logsin <= 24'd00186710;
                12'd1055: logsin <= 24'd00187067;
                12'd1056: logsin <= 24'd00187423;
                12'd1057: logsin <= 24'd00187780;
                12'd1058: logsin <= 24'd00188138;
                12'd1059: logsin <= 24'd00188495;
                12'd1060: logsin <= 24'd00188853;
                12'd1061: logsin <= 24'd00189212;
                12'd1062: logsin <= 24'd00189570;
                12'd1063: logsin <= 24'd00189930;
                12'd1064: logsin <= 24'd00190289;
                12'd1065: logsin <= 24'd00190649;
                12'd1066: logsin <= 24'd00191009;
                12'd1067: logsin <= 24'd00191369;
                12'd1068: logsin <= 24'd00191730;
                12'd1069: logsin <= 24'd00192091;
                12'd1070: logsin <= 24'd00192453;
                12'd1071: logsin <= 24'd00192814;
                12'd1072: logsin <= 24'd00193177;
                12'd1073: logsin <= 24'd00193539;
                12'd1074: logsin <= 24'd00193902;
                12'd1075: logsin <= 24'd00194265;
                12'd1076: logsin <= 24'd00194629;
                12'd1077: logsin <= 24'd00194993;
                12'd1078: logsin <= 24'd00195357;
                12'd1079: logsin <= 24'd00195721;
                12'd1080: logsin <= 24'd00196086;
                12'd1081: logsin <= 24'd00196452;
                12'd1082: logsin <= 24'd00196817;
                12'd1083: logsin <= 24'd00197183;
                12'd1084: logsin <= 24'd00197549;
                12'd1085: logsin <= 24'd00197916;
                12'd1086: logsin <= 24'd00198283;
                12'd1087: logsin <= 24'd00198650;
                12'd1088: logsin <= 24'd00199018;
                12'd1089: logsin <= 24'd00199386;
                12'd1090: logsin <= 24'd00199754;
                12'd1091: logsin <= 24'd00200123;
                12'd1092: logsin <= 24'd00200492;
                12'd1093: logsin <= 24'd00200862;
                12'd1094: logsin <= 24'd00201231;
                12'd1095: logsin <= 24'd00201601;
                12'd1096: logsin <= 24'd00201972;
                12'd1097: logsin <= 24'd00202343;
                12'd1098: logsin <= 24'd00202714;
                12'd1099: logsin <= 24'd00203085;
                12'd1100: logsin <= 24'd00203457;
                12'd1101: logsin <= 24'd00203829;
                12'd1102: logsin <= 24'd00204202;
                12'd1103: logsin <= 24'd00204575;
                12'd1104: logsin <= 24'd00204948;
                12'd1105: logsin <= 24'd00205321;
                12'd1106: logsin <= 24'd00205695;
                12'd1107: logsin <= 24'd00206069;
                12'd1108: logsin <= 24'd00206444;
                12'd1109: logsin <= 24'd00206819;
                12'd1110: logsin <= 24'd00207194;
                12'd1111: logsin <= 24'd00207570;
                12'd1112: logsin <= 24'd00207946;
                12'd1113: logsin <= 24'd00208322;
                12'd1114: logsin <= 24'd00208699;
                12'd1115: logsin <= 24'd00209076;
                12'd1116: logsin <= 24'd00209453;
                12'd1117: logsin <= 24'd00209831;
                12'd1118: logsin <= 24'd00210209;
                12'd1119: logsin <= 24'd00210587;
                12'd1120: logsin <= 24'd00210966;
                12'd1121: logsin <= 24'd00211345;
                12'd1122: logsin <= 24'd00211724;
                12'd1123: logsin <= 24'd00212104;
                12'd1124: logsin <= 24'd00212484;
                12'd1125: logsin <= 24'd00212865;
                12'd1126: logsin <= 24'd00213246;
                12'd1127: logsin <= 24'd00213627;
                12'd1128: logsin <= 24'd00214008;
                12'd1129: logsin <= 24'd00214390;
                12'd1130: logsin <= 24'd00214772;
                12'd1131: logsin <= 24'd00215155;
                12'd1132: logsin <= 24'd00215538;
                12'd1133: logsin <= 24'd00215921;
                12'd1134: logsin <= 24'd00216304;
                12'd1135: logsin <= 24'd00216688;
                12'd1136: logsin <= 24'd00217072;
                12'd1137: logsin <= 24'd00217457;
                12'd1138: logsin <= 24'd00217842;
                12'd1139: logsin <= 24'd00218227;
                12'd1140: logsin <= 24'd00218613;
                12'd1141: logsin <= 24'd00218999;
                12'd1142: logsin <= 24'd00219385;
                12'd1143: logsin <= 24'd00219772;
                12'd1144: logsin <= 24'd00220159;
                12'd1145: logsin <= 24'd00220546;
                12'd1146: logsin <= 24'd00220934;
                12'd1147: logsin <= 24'd00221322;
                12'd1148: logsin <= 24'd00221710;
                12'd1149: logsin <= 24'd00222099;
                12'd1150: logsin <= 24'd00222488;
                12'd1151: logsin <= 24'd00222878;
                12'd1152: logsin <= 24'd00223268;
                12'd1153: logsin <= 24'd00223658;
                12'd1154: logsin <= 24'd00224048;
                12'd1155: logsin <= 24'd00224439;
                12'd1156: logsin <= 24'd00224830;
                12'd1157: logsin <= 24'd00225222;
                12'd1158: logsin <= 24'd00225613;
                12'd1159: logsin <= 24'd00226006;
                12'd1160: logsin <= 24'd00226398;
                12'd1161: logsin <= 24'd00226791;
                12'd1162: logsin <= 24'd00227184;
                12'd1163: logsin <= 24'd00227578;
                12'd1164: logsin <= 24'd00227972;
                12'd1165: logsin <= 24'd00228366;
                12'd1166: logsin <= 24'd00228761;
                12'd1167: logsin <= 24'd00229156;
                12'd1168: logsin <= 24'd00229551;
                12'd1169: logsin <= 24'd00229947;
                12'd1170: logsin <= 24'd00230343;
                12'd1171: logsin <= 24'd00230739;
                12'd1172: logsin <= 24'd00231136;
                12'd1173: logsin <= 24'd00231533;
                12'd1174: logsin <= 24'd00231930;
                12'd1175: logsin <= 24'd00232328;
                12'd1176: logsin <= 24'd00232726;
                12'd1177: logsin <= 24'd00233124;
                12'd1178: logsin <= 24'd00233523;
                12'd1179: logsin <= 24'd00233922;
                12'd1180: logsin <= 24'd00234322;
                12'd1181: logsin <= 24'd00234722;
                12'd1182: logsin <= 24'd00235122;
                12'd1183: logsin <= 24'd00235522;
                12'd1184: logsin <= 24'd00235923;
                12'd1185: logsin <= 24'd00236324;
                12'd1186: logsin <= 24'd00236726;
                12'd1187: logsin <= 24'd00237128;
                12'd1188: logsin <= 24'd00237530;
                12'd1189: logsin <= 24'd00237933;
                12'd1190: logsin <= 24'd00238336;
                12'd1191: logsin <= 24'd00238739;
                12'd1192: logsin <= 24'd00239142;
                12'd1193: logsin <= 24'd00239546;
                12'd1194: logsin <= 24'd00239951;
                12'd1195: logsin <= 24'd00240355;
                12'd1196: logsin <= 24'd00240760;
                12'd1197: logsin <= 24'd00241166;
                12'd1198: logsin <= 24'd00241571;
                12'd1199: logsin <= 24'd00241978;
                12'd1200: logsin <= 24'd00242384;
                12'd1201: logsin <= 24'd00242791;
                12'd1202: logsin <= 24'd00243198;
                12'd1203: logsin <= 24'd00243605;
                12'd1204: logsin <= 24'd00244013;
                12'd1205: logsin <= 24'd00244421;
                12'd1206: logsin <= 24'd00244830;
                12'd1207: logsin <= 24'd00245238;
                12'd1208: logsin <= 24'd00245648;
                12'd1209: logsin <= 24'd00246057;
                12'd1210: logsin <= 24'd00246467;
                12'd1211: logsin <= 24'd00246877;
                12'd1212: logsin <= 24'd00247288;
                12'd1213: logsin <= 24'd00247699;
                12'd1214: logsin <= 24'd00248110;
                12'd1215: logsin <= 24'd00248521;
                12'd1216: logsin <= 24'd00248933;
                12'd1217: logsin <= 24'd00249346;
                12'd1218: logsin <= 24'd00249758;
                12'd1219: logsin <= 24'd00250171;
                12'd1220: logsin <= 24'd00250585;
                12'd1221: logsin <= 24'd00250998;
                12'd1222: logsin <= 24'd00251412;
                12'd1223: logsin <= 24'd00251827;
                12'd1224: logsin <= 24'd00252241;
                12'd1225: logsin <= 24'd00252656;
                12'd1226: logsin <= 24'd00253072;
                12'd1227: logsin <= 24'd00253487;
                12'd1228: logsin <= 24'd00253904;
                12'd1229: logsin <= 24'd00254320;
                12'd1230: logsin <= 24'd00254737;
                12'd1231: logsin <= 24'd00255154;
                12'd1232: logsin <= 24'd00255571;
                12'd1233: logsin <= 24'd00255989;
                12'd1234: logsin <= 24'd00256407;
                12'd1235: logsin <= 24'd00256826;
                12'd1236: logsin <= 24'd00257245;
                12'd1237: logsin <= 24'd00257664;
                12'd1238: logsin <= 24'd00258084;
                12'd1239: logsin <= 24'd00258503;
                12'd1240: logsin <= 24'd00258924;
                12'd1241: logsin <= 24'd00259344;
                12'd1242: logsin <= 24'd00259765;
                12'd1243: logsin <= 24'd00260187;
                12'd1244: logsin <= 24'd00260608;
                12'd1245: logsin <= 24'd00261030;
                12'd1246: logsin <= 24'd00261453;
                12'd1247: logsin <= 24'd00261875;
                12'd1248: logsin <= 24'd00262298;
                12'd1249: logsin <= 24'd00262722;
                12'd1250: logsin <= 24'd00263145;
                12'd1251: logsin <= 24'd00263569;
                12'd1252: logsin <= 24'd00263994;
                12'd1253: logsin <= 24'd00264419;
                12'd1254: logsin <= 24'd00264844;
                12'd1255: logsin <= 24'd00265269;
                12'd1256: logsin <= 24'd00265695;
                12'd1257: logsin <= 24'd00266121;
                12'd1258: logsin <= 24'd00266548;
                12'd1259: logsin <= 24'd00266974;
                12'd1260: logsin <= 24'd00267402;
                12'd1261: logsin <= 24'd00267829;
                12'd1262: logsin <= 24'd00268257;
                12'd1263: logsin <= 24'd00268685;
                12'd1264: logsin <= 24'd00269114;
                12'd1265: logsin <= 24'd00269543;
                12'd1266: logsin <= 24'd00269972;
                12'd1267: logsin <= 24'd00270402;
                12'd1268: logsin <= 24'd00270832;
                12'd1269: logsin <= 24'd00271262;
                12'd1270: logsin <= 24'd00271693;
                12'd1271: logsin <= 24'd00272124;
                12'd1272: logsin <= 24'd00272555;
                12'd1273: logsin <= 24'd00272987;
                12'd1274: logsin <= 24'd00273419;
                12'd1275: logsin <= 24'd00273851;
                12'd1276: logsin <= 24'd00274284;
                12'd1277: logsin <= 24'd00274717;
                12'd1278: logsin <= 24'd00275150;
                12'd1279: logsin <= 24'd00275584;
                12'd1280: logsin <= 24'd00276018;
                12'd1281: logsin <= 24'd00276453;
                12'd1282: logsin <= 24'd00276888;
                12'd1283: logsin <= 24'd00277323;
                12'd1284: logsin <= 24'd00277758;
                12'd1285: logsin <= 24'd00278194;
                12'd1286: logsin <= 24'd00278630;
                12'd1287: logsin <= 24'd00279067;
                12'd1288: logsin <= 24'd00279504;
                12'd1289: logsin <= 24'd00279941;
                12'd1290: logsin <= 24'd00280379;
                12'd1291: logsin <= 24'd00280817;
                12'd1292: logsin <= 24'd00281255;
                12'd1293: logsin <= 24'd00281694;
                12'd1294: logsin <= 24'd00282133;
                12'd1295: logsin <= 24'd00282572;
                12'd1296: logsin <= 24'd00283012;
                12'd1297: logsin <= 24'd00283452;
                12'd1298: logsin <= 24'd00283892;
                12'd1299: logsin <= 24'd00284333;
                12'd1300: logsin <= 24'd00284774;
                12'd1301: logsin <= 24'd00285215;
                12'd1302: logsin <= 24'd00285657;
                12'd1303: logsin <= 24'd00286099;
                12'd1304: logsin <= 24'd00286542;
                12'd1305: logsin <= 24'd00286984;
                12'd1306: logsin <= 24'd00287428;
                12'd1307: logsin <= 24'd00287871;
                12'd1308: logsin <= 24'd00288315;
                12'd1309: logsin <= 24'd00288759;
                12'd1310: logsin <= 24'd00289204;
                12'd1311: logsin <= 24'd00289649;
                12'd1312: logsin <= 24'd00290094;
                12'd1313: logsin <= 24'd00290539;
                12'd1314: logsin <= 24'd00290985;
                12'd1315: logsin <= 24'd00291432;
                12'd1316: logsin <= 24'd00291878;
                12'd1317: logsin <= 24'd00292325;
                12'd1318: logsin <= 24'd00292773;
                12'd1319: logsin <= 24'd00293220;
                12'd1320: logsin <= 24'd00293668;
                12'd1321: logsin <= 24'd00294117;
                12'd1322: logsin <= 24'd00294565;
                12'd1323: logsin <= 24'd00295014;
                12'd1324: logsin <= 24'd00295464;
                12'd1325: logsin <= 24'd00295914;
                12'd1326: logsin <= 24'd00296364;
                12'd1327: logsin <= 24'd00296814;
                12'd1328: logsin <= 24'd00297265;
                12'd1329: logsin <= 24'd00297716;
                12'd1330: logsin <= 24'd00298168;
                12'd1331: logsin <= 24'd00298619;
                12'd1332: logsin <= 24'd00299072;
                12'd1333: logsin <= 24'd00299524;
                12'd1334: logsin <= 24'd00299977;
                12'd1335: logsin <= 24'd00300430;
                12'd1336: logsin <= 24'd00300884;
                12'd1337: logsin <= 24'd00301338;
                12'd1338: logsin <= 24'd00301792;
                12'd1339: logsin <= 24'd00302247;
                12'd1340: logsin <= 24'd00302702;
                12'd1341: logsin <= 24'd00303157;
                12'd1342: logsin <= 24'd00303613;
                12'd1343: logsin <= 24'd00304069;
                12'd1344: logsin <= 24'd00304525;
                12'd1345: logsin <= 24'd00304982;
                12'd1346: logsin <= 24'd00305439;
                12'd1347: logsin <= 24'd00305896;
                12'd1348: logsin <= 24'd00306354;
                12'd1349: logsin <= 24'd00306812;
                12'd1350: logsin <= 24'd00307270;
                12'd1351: logsin <= 24'd00307729;
                12'd1352: logsin <= 24'd00308188;
                12'd1353: logsin <= 24'd00308648;
                12'd1354: logsin <= 24'd00309108;
                12'd1355: logsin <= 24'd00309568;
                12'd1356: logsin <= 24'd00310028;
                12'd1357: logsin <= 24'd00310489;
                12'd1358: logsin <= 24'd00310950;
                12'd1359: logsin <= 24'd00311412;
                12'd1360: logsin <= 24'd00311874;
                12'd1361: logsin <= 24'd00312336;
                12'd1362: logsin <= 24'd00312799;
                12'd1363: logsin <= 24'd00313262;
                12'd1364: logsin <= 24'd00313725;
                12'd1365: logsin <= 24'd00314189;
                12'd1366: logsin <= 24'd00314653;
                12'd1367: logsin <= 24'd00315117;
                12'd1368: logsin <= 24'd00315582;
                12'd1369: logsin <= 24'd00316047;
                12'd1370: logsin <= 24'd00316512;
                12'd1371: logsin <= 24'd00316978;
                12'd1372: logsin <= 24'd00317444;
                12'd1373: logsin <= 24'd00317910;
                12'd1374: logsin <= 24'd00318377;
                12'd1375: logsin <= 24'd00318844;
                12'd1376: logsin <= 24'd00319312;
                12'd1377: logsin <= 24'd00319780;
                12'd1378: logsin <= 24'd00320248;
                12'd1379: logsin <= 24'd00320716;
                12'd1380: logsin <= 24'd00321185;
                12'd1381: logsin <= 24'd00321654;
                12'd1382: logsin <= 24'd00322124;
                12'd1383: logsin <= 24'd00322594;
                12'd1384: logsin <= 24'd00323064;
                12'd1385: logsin <= 24'd00323535;
                12'd1386: logsin <= 24'd00324006;
                12'd1387: logsin <= 24'd00324477;
                12'd1388: logsin <= 24'd00324949;
                12'd1389: logsin <= 24'd00325421;
                12'd1390: logsin <= 24'd00325893;
                12'd1391: logsin <= 24'd00326366;
                12'd1392: logsin <= 24'd00326839;
                12'd1393: logsin <= 24'd00327312;
                12'd1394: logsin <= 24'd00327786;
                12'd1395: logsin <= 24'd00328260;
                12'd1396: logsin <= 24'd00328734;
                12'd1397: logsin <= 24'd00329209;
                12'd1398: logsin <= 24'd00329684;
                12'd1399: logsin <= 24'd00330160;
                12'd1400: logsin <= 24'd00330636;
                12'd1401: logsin <= 24'd00331112;
                12'd1402: logsin <= 24'd00331588;
                12'd1403: logsin <= 24'd00332065;
                12'd1404: logsin <= 24'd00332542;
                12'd1405: logsin <= 24'd00333020;
                12'd1406: logsin <= 24'd00333498;
                12'd1407: logsin <= 24'd00333976;
                12'd1408: logsin <= 24'd00334455;
                12'd1409: logsin <= 24'd00334934;
                12'd1410: logsin <= 24'd00335413;
                12'd1411: logsin <= 24'd00335893;
                12'd1412: logsin <= 24'd00336372;
                12'd1413: logsin <= 24'd00336853;
                12'd1414: logsin <= 24'd00337334;
                12'd1415: logsin <= 24'd00337815;
                12'd1416: logsin <= 24'd00338296;
                12'd1417: logsin <= 24'd00338778;
                12'd1418: logsin <= 24'd00339260;
                12'd1419: logsin <= 24'd00339742;
                12'd1420: logsin <= 24'd00340225;
                12'd1421: logsin <= 24'd00340708;
                12'd1422: logsin <= 24'd00341192;
                12'd1423: logsin <= 24'd00341675;
                12'd1424: logsin <= 24'd00342160;
                12'd1425: logsin <= 24'd00342644;
                12'd1426: logsin <= 24'd00343129;
                12'd1427: logsin <= 24'd00343614;
                12'd1428: logsin <= 24'd00344100;
                12'd1429: logsin <= 24'd00344586;
                12'd1430: logsin <= 24'd00345072;
                12'd1431: logsin <= 24'd00345558;
                12'd1432: logsin <= 24'd00346045;
                12'd1433: logsin <= 24'd00346533;
                12'd1434: logsin <= 24'd00347020;
                12'd1435: logsin <= 24'd00347508;
                12'd1436: logsin <= 24'd00347997;
                12'd1437: logsin <= 24'd00348485;
                12'd1438: logsin <= 24'd00348974;
                12'd1439: logsin <= 24'd00349464;
                12'd1440: logsin <= 24'd00349953;
                12'd1441: logsin <= 24'd00350443;
                12'd1442: logsin <= 24'd00350934;
                12'd1443: logsin <= 24'd00351425;
                12'd1444: logsin <= 24'd00351916;
                12'd1445: logsin <= 24'd00352407;
                12'd1446: logsin <= 24'd00352899;
                12'd1447: logsin <= 24'd00353391;
                12'd1448: logsin <= 24'd00353884;
                12'd1449: logsin <= 24'd00354377;
                12'd1450: logsin <= 24'd00354870;
                12'd1451: logsin <= 24'd00355363;
                12'd1452: logsin <= 24'd00355857;
                12'd1453: logsin <= 24'd00356351;
                12'd1454: logsin <= 24'd00356846;
                12'd1455: logsin <= 24'd00357341;
                12'd1456: logsin <= 24'd00357836;
                12'd1457: logsin <= 24'd00358332;
                12'd1458: logsin <= 24'd00358828;
                12'd1459: logsin <= 24'd00359324;
                12'd1460: logsin <= 24'd00359821;
                12'd1461: logsin <= 24'd00360318;
                12'd1462: logsin <= 24'd00360815;
                12'd1463: logsin <= 24'd00361313;
                12'd1464: logsin <= 24'd00361811;
                12'd1465: logsin <= 24'd00362309;
                12'd1466: logsin <= 24'd00362808;
                12'd1467: logsin <= 24'd00363307;
                12'd1468: logsin <= 24'd00363807;
                12'd1469: logsin <= 24'd00364307;
                12'd1470: logsin <= 24'd00364807;
                12'd1471: logsin <= 24'd00365307;
                12'd1472: logsin <= 24'd00365808;
                12'd1473: logsin <= 24'd00366309;
                12'd1474: logsin <= 24'd00366811;
                12'd1475: logsin <= 24'd00367313;
                12'd1476: logsin <= 24'd00367815;
                12'd1477: logsin <= 24'd00368318;
                12'd1478: logsin <= 24'd00368820;
                12'd1479: logsin <= 24'd00369324;
                12'd1480: logsin <= 24'd00369827;
                12'd1481: logsin <= 24'd00370331;
                12'd1482: logsin <= 24'd00370836;
                12'd1483: logsin <= 24'd00371340;
                12'd1484: logsin <= 24'd00371845;
                12'd1485: logsin <= 24'd00372351;
                12'd1486: logsin <= 24'd00372856;
                12'd1487: logsin <= 24'd00373363;
                12'd1488: logsin <= 24'd00373869;
                12'd1489: logsin <= 24'd00374376;
                12'd1490: logsin <= 24'd00374883;
                12'd1491: logsin <= 24'd00375390;
                12'd1492: logsin <= 24'd00375898;
                12'd1493: logsin <= 24'd00376406;
                12'd1494: logsin <= 24'd00376915;
                12'd1495: logsin <= 24'd00377423;
                12'd1496: logsin <= 24'd00377933;
                12'd1497: logsin <= 24'd00378442;
                12'd1498: logsin <= 24'd00378952;
                12'd1499: logsin <= 24'd00379462;
                12'd1500: logsin <= 24'd00379973;
                12'd1501: logsin <= 24'd00380484;
                12'd1502: logsin <= 24'd00380995;
                12'd1503: logsin <= 24'd00381507;
                12'd1504: logsin <= 24'd00382019;
                12'd1505: logsin <= 24'd00382531;
                12'd1506: logsin <= 24'd00383044;
                12'd1507: logsin <= 24'd00383557;
                12'd1508: logsin <= 24'd00384070;
                12'd1509: logsin <= 24'd00384584;
                12'd1510: logsin <= 24'd00385098;
                12'd1511: logsin <= 24'd00385612;
                12'd1512: logsin <= 24'd00386127;
                12'd1513: logsin <= 24'd00386642;
                12'd1514: logsin <= 24'd00387157;
                12'd1515: logsin <= 24'd00387673;
                12'd1516: logsin <= 24'd00388189;
                12'd1517: logsin <= 24'd00388706;
                12'd1518: logsin <= 24'd00389223;
                12'd1519: logsin <= 24'd00389740;
                12'd1520: logsin <= 24'd00390257;
                12'd1521: logsin <= 24'd00390775;
                12'd1522: logsin <= 24'd00391293;
                12'd1523: logsin <= 24'd00391812;
                12'd1524: logsin <= 24'd00392331;
                12'd1525: logsin <= 24'd00392850;
                12'd1526: logsin <= 24'd00393370;
                12'd1527: logsin <= 24'd00393890;
                12'd1528: logsin <= 24'd00394410;
                12'd1529: logsin <= 24'd00394931;
                12'd1530: logsin <= 24'd00395452;
                12'd1531: logsin <= 24'd00395973;
                12'd1532: logsin <= 24'd00396495;
                12'd1533: logsin <= 24'd00397017;
                12'd1534: logsin <= 24'd00397539;
                12'd1535: logsin <= 24'd00398062;
                12'd1536: logsin <= 24'd00398585;
                12'd1537: logsin <= 24'd00399108;
                12'd1538: logsin <= 24'd00399632;
                12'd1539: logsin <= 24'd00400156;
                12'd1540: logsin <= 24'd00400681;
                12'd1541: logsin <= 24'd00401205;
                12'd1542: logsin <= 24'd00401731;
                12'd1543: logsin <= 24'd00402256;
                12'd1544: logsin <= 24'd00402782;
                12'd1545: logsin <= 24'd00403308;
                12'd1546: logsin <= 24'd00403835;
                12'd1547: logsin <= 24'd00404362;
                12'd1548: logsin <= 24'd00404889;
                12'd1549: logsin <= 24'd00405416;
                12'd1550: logsin <= 24'd00405944;
                12'd1551: logsin <= 24'd00406473;
                12'd1552: logsin <= 24'd00407001;
                12'd1553: logsin <= 24'd00407530;
                12'd1554: logsin <= 24'd00408060;
                12'd1555: logsin <= 24'd00408589;
                12'd1556: logsin <= 24'd00409119;
                12'd1557: logsin <= 24'd00409650;
                12'd1558: logsin <= 24'd00410180;
                12'd1559: logsin <= 24'd00410711;
                12'd1560: logsin <= 24'd00411243;
                12'd1561: logsin <= 24'd00411774;
                12'd1562: logsin <= 24'd00412307;
                12'd1563: logsin <= 24'd00412839;
                12'd1564: logsin <= 24'd00413372;
                12'd1565: logsin <= 24'd00413905;
                12'd1566: logsin <= 24'd00414438;
                12'd1567: logsin <= 24'd00414972;
                12'd1568: logsin <= 24'd00415506;
                12'd1569: logsin <= 24'd00416041;
                12'd1570: logsin <= 24'd00416576;
                12'd1571: logsin <= 24'd00417111;
                12'd1572: logsin <= 24'd00417647;
                12'd1573: logsin <= 24'd00418182;
                12'd1574: logsin <= 24'd00418719;
                12'd1575: logsin <= 24'd00419255;
                12'd1576: logsin <= 24'd00419792;
                12'd1577: logsin <= 24'd00420330;
                12'd1578: logsin <= 24'd00420867;
                12'd1579: logsin <= 24'd00421405;
                12'd1580: logsin <= 24'd00421944;
                12'd1581: logsin <= 24'd00422482;
                12'd1582: logsin <= 24'd00423021;
                12'd1583: logsin <= 24'd00423561;
                12'd1584: logsin <= 24'd00424100;
                12'd1585: logsin <= 24'd00424640;
                12'd1586: logsin <= 24'd00425181;
                12'd1587: logsin <= 24'd00425722;
                12'd1588: logsin <= 24'd00426263;
                12'd1589: logsin <= 24'd00426804;
                12'd1590: logsin <= 24'd00427346;
                12'd1591: logsin <= 24'd00427888;
                12'd1592: logsin <= 24'd00428431;
                12'd1593: logsin <= 24'd00428973;
                12'd1594: logsin <= 24'd00429517;
                12'd1595: logsin <= 24'd00430060;
                12'd1596: logsin <= 24'd00430604;
                12'd1597: logsin <= 24'd00431148;
                12'd1598: logsin <= 24'd00431693;
                12'd1599: logsin <= 24'd00432238;
                12'd1600: logsin <= 24'd00432783;
                12'd1601: logsin <= 24'd00433329;
                12'd1602: logsin <= 24'd00433875;
                12'd1603: logsin <= 24'd00434421;
                12'd1604: logsin <= 24'd00434967;
                12'd1605: logsin <= 24'd00435514;
                12'd1606: logsin <= 24'd00436062;
                12'd1607: logsin <= 24'd00436609;
                12'd1608: logsin <= 24'd00437157;
                12'd1609: logsin <= 24'd00437706;
                12'd1610: logsin <= 24'd00438255;
                12'd1611: logsin <= 24'd00438804;
                12'd1612: logsin <= 24'd00439353;
                12'd1613: logsin <= 24'd00439903;
                12'd1614: logsin <= 24'd00440453;
                12'd1615: logsin <= 24'd00441003;
                12'd1616: logsin <= 24'd00441554;
                12'd1617: logsin <= 24'd00442105;
                12'd1618: logsin <= 24'd00442657;
                12'd1619: logsin <= 24'd00443209;
                12'd1620: logsin <= 24'd00443761;
                12'd1621: logsin <= 24'd00444313;
                12'd1622: logsin <= 24'd00444866;
                12'd1623: logsin <= 24'd00445419;
                12'd1624: logsin <= 24'd00445973;
                12'd1625: logsin <= 24'd00446527;
                12'd1626: logsin <= 24'd00447081;
                12'd1627: logsin <= 24'd00447636;
                12'd1628: logsin <= 24'd00448191;
                12'd1629: logsin <= 24'd00448746;
                12'd1630: logsin <= 24'd00449302;
                12'd1631: logsin <= 24'd00449858;
                12'd1632: logsin <= 24'd00450414;
                12'd1633: logsin <= 24'd00450971;
                12'd1634: logsin <= 24'd00451528;
                12'd1635: logsin <= 24'd00452085;
                12'd1636: logsin <= 24'd00452643;
                12'd1637: logsin <= 24'd00453201;
                12'd1638: logsin <= 24'd00453759;
                12'd1639: logsin <= 24'd00454318;
                12'd1640: logsin <= 24'd00454877;
                12'd1641: logsin <= 24'd00455436;
                12'd1642: logsin <= 24'd00455996;
                12'd1643: logsin <= 24'd00456556;
                12'd1644: logsin <= 24'd00457117;
                12'd1645: logsin <= 24'd00457678;
                12'd1646: logsin <= 24'd00458239;
                12'd1647: logsin <= 24'd00458800;
                12'd1648: logsin <= 24'd00459362;
                12'd1649: logsin <= 24'd00459924;
                12'd1650: logsin <= 24'd00460487;
                12'd1651: logsin <= 24'd00461050;
                12'd1652: logsin <= 24'd00461613;
                12'd1653: logsin <= 24'd00462177;
                12'd1654: logsin <= 24'd00462741;
                12'd1655: logsin <= 24'd00463305;
                12'd1656: logsin <= 24'd00463869;
                12'd1657: logsin <= 24'd00464434;
                12'd1658: logsin <= 24'd00465000;
                12'd1659: logsin <= 24'd00465565;
                12'd1660: logsin <= 24'd00466131;
                12'd1661: logsin <= 24'd00466698;
                12'd1662: logsin <= 24'd00467264;
                12'd1663: logsin <= 24'd00467831;
                12'd1664: logsin <= 24'd00468399;
                12'd1665: logsin <= 24'd00468966;
                12'd1666: logsin <= 24'd00469535;
                12'd1667: logsin <= 24'd00470103;
                12'd1668: logsin <= 24'd00470672;
                12'd1669: logsin <= 24'd00471241;
                12'd1670: logsin <= 24'd00471810;
                12'd1671: logsin <= 24'd00472380;
                12'd1672: logsin <= 24'd00472950;
                12'd1673: logsin <= 24'd00473521;
                12'd1674: logsin <= 24'd00474091;
                12'd1675: logsin <= 24'd00474663;
                12'd1676: logsin <= 24'd00475234;
                12'd1677: logsin <= 24'd00475806;
                12'd1678: logsin <= 24'd00476378;
                12'd1679: logsin <= 24'd00476951;
                12'd1680: logsin <= 24'd00477524;
                12'd1681: logsin <= 24'd00478097;
                12'd1682: logsin <= 24'd00478670;
                12'd1683: logsin <= 24'd00479244;
                12'd1684: logsin <= 24'd00479819;
                12'd1685: logsin <= 24'd00480393;
                12'd1686: logsin <= 24'd00480968;
                12'd1687: logsin <= 24'd00481543;
                12'd1688: logsin <= 24'd00482119;
                12'd1689: logsin <= 24'd00482695;
                12'd1690: logsin <= 24'd00483271;
                12'd1691: logsin <= 24'd00483848;
                12'd1692: logsin <= 24'd00484425;
                12'd1693: logsin <= 24'd00485002;
                12'd1694: logsin <= 24'd00485580;
                12'd1695: logsin <= 24'd00486158;
                12'd1696: logsin <= 24'd00486737;
                12'd1697: logsin <= 24'd00487315;
                12'd1698: logsin <= 24'd00487894;
                12'd1699: logsin <= 24'd00488474;
                12'd1700: logsin <= 24'd00489054;
                12'd1701: logsin <= 24'd00489634;
                12'd1702: logsin <= 24'd00490214;
                12'd1703: logsin <= 24'd00490795;
                12'd1704: logsin <= 24'd00491376;
                12'd1705: logsin <= 24'd00491958;
                12'd1706: logsin <= 24'd00492539;
                12'd1707: logsin <= 24'd00493122;
                12'd1708: logsin <= 24'd00493704;
                12'd1709: logsin <= 24'd00494287;
                12'd1710: logsin <= 24'd00494870;
                12'd1711: logsin <= 24'd00495454;
                12'd1712: logsin <= 24'd00496038;
                12'd1713: logsin <= 24'd00496622;
                12'd1714: logsin <= 24'd00497206;
                12'd1715: logsin <= 24'd00497791;
                12'd1716: logsin <= 24'd00498377;
                12'd1717: logsin <= 24'd00498962;
                12'd1718: logsin <= 24'd00499548;
                12'd1719: logsin <= 24'd00500135;
                12'd1720: logsin <= 24'd00500721;
                12'd1721: logsin <= 24'd00501308;
                12'd1722: logsin <= 24'd00501895;
                12'd1723: logsin <= 24'd00502483;
                12'd1724: logsin <= 24'd00503071;
                12'd1725: logsin <= 24'd00503659;
                12'd1726: logsin <= 24'd00504248;
                12'd1727: logsin <= 24'd00504837;
                12'd1728: logsin <= 24'd00505427;
                12'd1729: logsin <= 24'd00506016;
                12'd1730: logsin <= 24'd00506606;
                12'd1731: logsin <= 24'd00507197;
                12'd1732: logsin <= 24'd00507788;
                12'd1733: logsin <= 24'd00508379;
                12'd1734: logsin <= 24'd00508970;
                12'd1735: logsin <= 24'd00509562;
                12'd1736: logsin <= 24'd00510154;
                12'd1737: logsin <= 24'd00510746;
                12'd1738: logsin <= 24'd00511339;
                12'd1739: logsin <= 24'd00511932;
                12'd1740: logsin <= 24'd00512526;
                12'd1741: logsin <= 24'd00513120;
                12'd1742: logsin <= 24'd00513714;
                12'd1743: logsin <= 24'd00514308;
                12'd1744: logsin <= 24'd00514903;
                12'd1745: logsin <= 24'd00515499;
                12'd1746: logsin <= 24'd00516094;
                12'd1747: logsin <= 24'd00516690;
                12'd1748: logsin <= 24'd00517286;
                12'd1749: logsin <= 24'd00517883;
                12'd1750: logsin <= 24'd00518480;
                12'd1751: logsin <= 24'd00519077;
                12'd1752: logsin <= 24'd00519675;
                12'd1753: logsin <= 24'd00520272;
                12'd1754: logsin <= 24'd00520871;
                12'd1755: logsin <= 24'd00521469;
                12'd1756: logsin <= 24'd00522068;
                12'd1757: logsin <= 24'd00522668;
                12'd1758: logsin <= 24'd00523267;
                12'd1759: logsin <= 24'd00523867;
                12'd1760: logsin <= 24'd00524468;
                12'd1761: logsin <= 24'd00525068;
                12'd1762: logsin <= 24'd00525669;
                12'd1763: logsin <= 24'd00526271;
                12'd1764: logsin <= 24'd00526872;
                12'd1765: logsin <= 24'd00527474;
                12'd1766: logsin <= 24'd00528077;
                12'd1767: logsin <= 24'd00528680;
                12'd1768: logsin <= 24'd00529283;
                12'd1769: logsin <= 24'd00529886;
                12'd1770: logsin <= 24'd00530490;
                12'd1771: logsin <= 24'd00531094;
                12'd1772: logsin <= 24'd00531698;
                12'd1773: logsin <= 24'd00532303;
                12'd1774: logsin <= 24'd00532908;
                12'd1775: logsin <= 24'd00533514;
                12'd1776: logsin <= 24'd00534119;
                12'd1777: logsin <= 24'd00534726;
                12'd1778: logsin <= 24'd00535332;
                12'd1779: logsin <= 24'd00535939;
                12'd1780: logsin <= 24'd00536546;
                12'd1781: logsin <= 24'd00537154;
                12'd1782: logsin <= 24'd00537761;
                12'd1783: logsin <= 24'd00538370;
                12'd1784: logsin <= 24'd00538978;
                12'd1785: logsin <= 24'd00539587;
                12'd1786: logsin <= 24'd00540196;
                12'd1787: logsin <= 24'd00540806;
                12'd1788: logsin <= 24'd00541416;
                12'd1789: logsin <= 24'd00542026;
                12'd1790: logsin <= 24'd00542636;
                12'd1791: logsin <= 24'd00543247;
                12'd1792: logsin <= 24'd00543859;
                12'd1793: logsin <= 24'd00544470;
                12'd1794: logsin <= 24'd00545082;
                12'd1795: logsin <= 24'd00545694;
                12'd1796: logsin <= 24'd00546307;
                12'd1797: logsin <= 24'd00546920;
                12'd1798: logsin <= 24'd00547533;
                12'd1799: logsin <= 24'd00548147;
                12'd1800: logsin <= 24'd00548761;
                12'd1801: logsin <= 24'd00549375;
                12'd1802: logsin <= 24'd00549990;
                12'd1803: logsin <= 24'd00550605;
                12'd1804: logsin <= 24'd00551220;
                12'd1805: logsin <= 24'd00551836;
                12'd1806: logsin <= 24'd00552452;
                12'd1807: logsin <= 24'd00553068;
                12'd1808: logsin <= 24'd00553685;
                12'd1809: logsin <= 24'd00554302;
                12'd1810: logsin <= 24'd00554919;
                12'd1811: logsin <= 24'd00555537;
                12'd1812: logsin <= 24'd00556155;
                12'd1813: logsin <= 24'd00556773;
                12'd1814: logsin <= 24'd00557392;
                12'd1815: logsin <= 24'd00558011;
                12'd1816: logsin <= 24'd00558630;
                12'd1817: logsin <= 24'd00559250;
                12'd1818: logsin <= 24'd00559870;
                12'd1819: logsin <= 24'd00560491;
                12'd1820: logsin <= 24'd00561111;
                12'd1821: logsin <= 24'd00561732;
                12'd1822: logsin <= 24'd00562354;
                12'd1823: logsin <= 24'd00562976;
                12'd1824: logsin <= 24'd00563598;
                12'd1825: logsin <= 24'd00564220;
                12'd1826: logsin <= 24'd00564843;
                12'd1827: logsin <= 24'd00565466;
                12'd1828: logsin <= 24'd00566090;
                12'd1829: logsin <= 24'd00566713;
                12'd1830: logsin <= 24'd00567337;
                12'd1831: logsin <= 24'd00567962;
                12'd1832: logsin <= 24'd00568587;
                12'd1833: logsin <= 24'd00569212;
                12'd1834: logsin <= 24'd00569837;
                12'd1835: logsin <= 24'd00570463;
                12'd1836: logsin <= 24'd00571089;
                12'd1837: logsin <= 24'd00571716;
                12'd1838: logsin <= 24'd00572343;
                12'd1839: logsin <= 24'd00572970;
                12'd1840: logsin <= 24'd00573597;
                12'd1841: logsin <= 24'd00574225;
                12'd1842: logsin <= 24'd00574853;
                12'd1843: logsin <= 24'd00575482;
                12'd1844: logsin <= 24'd00576111;
                12'd1845: logsin <= 24'd00576740;
                12'd1846: logsin <= 24'd00577370;
                12'd1847: logsin <= 24'd00578000;
                12'd1848: logsin <= 24'd00578630;
                12'd1849: logsin <= 24'd00579260;
                12'd1850: logsin <= 24'd00579891;
                12'd1851: logsin <= 24'd00580522;
                12'd1852: logsin <= 24'd00581154;
                12'd1853: logsin <= 24'd00581786;
                12'd1854: logsin <= 24'd00582418;
                12'd1855: logsin <= 24'd00583051;
                12'd1856: logsin <= 24'd00583684;
                12'd1857: logsin <= 24'd00584317;
                12'd1858: logsin <= 24'd00584950;
                12'd1859: logsin <= 24'd00585584;
                12'd1860: logsin <= 24'd00586219;
                12'd1861: logsin <= 24'd00586853;
                12'd1862: logsin <= 24'd00587488;
                12'd1863: logsin <= 24'd00588123;
                12'd1864: logsin <= 24'd00588759;
                12'd1865: logsin <= 24'd00589395;
                12'd1866: logsin <= 24'd00590031;
                12'd1867: logsin <= 24'd00590668;
                12'd1868: logsin <= 24'd00591305;
                12'd1869: logsin <= 24'd00591942;
                12'd1870: logsin <= 24'd00592580;
                12'd1871: logsin <= 24'd00593218;
                12'd1872: logsin <= 24'd00593856;
                12'd1873: logsin <= 24'd00594495;
                12'd1874: logsin <= 24'd00595134;
                12'd1875: logsin <= 24'd00595773;
                12'd1876: logsin <= 24'd00596413;
                12'd1877: logsin <= 24'd00597053;
                12'd1878: logsin <= 24'd00597693;
                12'd1879: logsin <= 24'd00598333;
                12'd1880: logsin <= 24'd00598974;
                12'd1881: logsin <= 24'd00599616;
                12'd1882: logsin <= 24'd00600257;
                12'd1883: logsin <= 24'd00600899;
                12'd1884: logsin <= 24'd00601542;
                12'd1885: logsin <= 24'd00602184;
                12'd1886: logsin <= 24'd00602827;
                12'd1887: logsin <= 24'd00603471;
                12'd1888: logsin <= 24'd00604114;
                12'd1889: logsin <= 24'd00604758;
                12'd1890: logsin <= 24'd00605403;
                12'd1891: logsin <= 24'd00606047;
                12'd1892: logsin <= 24'd00606692;
                12'd1893: logsin <= 24'd00607338;
                12'd1894: logsin <= 24'd00607983;
                12'd1895: logsin <= 24'd00608629;
                12'd1896: logsin <= 24'd00609276;
                12'd1897: logsin <= 24'd00609922;
                12'd1898: logsin <= 24'd00610569;
                12'd1899: logsin <= 24'd00611217;
                12'd1900: logsin <= 24'd00611864;
                12'd1901: logsin <= 24'd00612512;
                12'd1902: logsin <= 24'd00613161;
                12'd1903: logsin <= 24'd00613809;
                12'd1904: logsin <= 24'd00614458;
                12'd1905: logsin <= 24'd00615108;
                12'd1906: logsin <= 24'd00615757;
                12'd1907: logsin <= 24'd00616407;
                12'd1908: logsin <= 24'd00617058;
                12'd1909: logsin <= 24'd00617708;
                12'd1910: logsin <= 24'd00618359;
                12'd1911: logsin <= 24'd00619011;
                12'd1912: logsin <= 24'd00619662;
                12'd1913: logsin <= 24'd00620314;
                12'd1914: logsin <= 24'd00620967;
                12'd1915: logsin <= 24'd00621619;
                12'd1916: logsin <= 24'd00622273;
                12'd1917: logsin <= 24'd00622926;
                12'd1918: logsin <= 24'd00623580;
                12'd1919: logsin <= 24'd00624234;
                12'd1920: logsin <= 24'd00624888;
                12'd1921: logsin <= 24'd00625543;
                12'd1922: logsin <= 24'd00626198;
                12'd1923: logsin <= 24'd00626853;
                12'd1924: logsin <= 24'd00627509;
                12'd1925: logsin <= 24'd00628165;
                12'd1926: logsin <= 24'd00628821;
                12'd1927: logsin <= 24'd00629478;
                12'd1928: logsin <= 24'd00630135;
                12'd1929: logsin <= 24'd00630792;
                12'd1930: logsin <= 24'd00631449;
                12'd1931: logsin <= 24'd00632107;
                12'd1932: logsin <= 24'd00632766;
                12'd1933: logsin <= 24'd00633424;
                12'd1934: logsin <= 24'd00634083;
                12'd1935: logsin <= 24'd00634743;
                12'd1936: logsin <= 24'd00635402;
                12'd1937: logsin <= 24'd00636062;
                12'd1938: logsin <= 24'd00636723;
                12'd1939: logsin <= 24'd00637383;
                12'd1940: logsin <= 24'd00638044;
                12'd1941: logsin <= 24'd00638706;
                12'd1942: logsin <= 24'd00639367;
                12'd1943: logsin <= 24'd00640029;
                12'd1944: logsin <= 24'd00640691;
                12'd1945: logsin <= 24'd00641354;
                12'd1946: logsin <= 24'd00642017;
                12'd1947: logsin <= 24'd00642680;
                12'd1948: logsin <= 24'd00643344;
                12'd1949: logsin <= 24'd00644008;
                12'd1950: logsin <= 24'd00644672;
                12'd1951: logsin <= 24'd00645337;
                12'd1952: logsin <= 24'd00646002;
                12'd1953: logsin <= 24'd00646667;
                12'd1954: logsin <= 24'd00647333;
                12'd1955: logsin <= 24'd00647999;
                12'd1956: logsin <= 24'd00648665;
                12'd1957: logsin <= 24'd00649331;
                12'd1958: logsin <= 24'd00649998;
                12'd1959: logsin <= 24'd00650665;
                12'd1960: logsin <= 24'd00651333;
                12'd1961: logsin <= 24'd00652001;
                12'd1962: logsin <= 24'd00652669;
                12'd1963: logsin <= 24'd00653338;
                12'd1964: logsin <= 24'd00654007;
                12'd1965: logsin <= 24'd00654676;
                12'd1966: logsin <= 24'd00655345;
                12'd1967: logsin <= 24'd00656015;
                12'd1968: logsin <= 24'd00656685;
                12'd1969: logsin <= 24'd00657356;
                12'd1970: logsin <= 24'd00658027;
                12'd1971: logsin <= 24'd00658698;
                12'd1972: logsin <= 24'd00659370;
                12'd1973: logsin <= 24'd00660041;
                12'd1974: logsin <= 24'd00660714;
                12'd1975: logsin <= 24'd00661386;
                12'd1976: logsin <= 24'd00662059;
                12'd1977: logsin <= 24'd00662732;
                12'd1978: logsin <= 24'd00663406;
                12'd1979: logsin <= 24'd00664079;
                12'd1980: logsin <= 24'd00664753;
                12'd1981: logsin <= 24'd00665428;
                12'd1982: logsin <= 24'd00666103;
                12'd1983: logsin <= 24'd00666778;
                12'd1984: logsin <= 24'd00667453;
                12'd1985: logsin <= 24'd00668129;
                12'd1986: logsin <= 24'd00668805;
                12'd1987: logsin <= 24'd00669482;
                12'd1988: logsin <= 24'd00670158;
                12'd1989: logsin <= 24'd00670835;
                12'd1990: logsin <= 24'd00671513;
                12'd1991: logsin <= 24'd00672191;
                12'd1992: logsin <= 24'd00672869;
                12'd1993: logsin <= 24'd00673547;
                12'd1994: logsin <= 24'd00674226;
                12'd1995: logsin <= 24'd00674905;
                12'd1996: logsin <= 24'd00675584;
                12'd1997: logsin <= 24'd00676264;
                12'd1998: logsin <= 24'd00676944;
                12'd1999: logsin <= 24'd00677624;
                12'd2000: logsin <= 24'd00678305;
                12'd2001: logsin <= 24'd00678986;
                12'd2002: logsin <= 24'd00679667;
                12'd2003: logsin <= 24'd00680349;
                12'd2004: logsin <= 24'd00681031;
                12'd2005: logsin <= 24'd00681713;
                12'd2006: logsin <= 24'd00682396;
                12'd2007: logsin <= 24'd00683079;
                12'd2008: logsin <= 24'd00683762;
                12'd2009: logsin <= 24'd00684445;
                12'd2010: logsin <= 24'd00685129;
                12'd2011: logsin <= 24'd00685814;
                12'd2012: logsin <= 24'd00686498;
                12'd2013: logsin <= 24'd00687183;
                12'd2014: logsin <= 24'd00687868;
                12'd2015: logsin <= 24'd00688554;
                12'd2016: logsin <= 24'd00689240;
                12'd2017: logsin <= 24'd00689926;
                12'd2018: logsin <= 24'd00690612;
                12'd2019: logsin <= 24'd00691299;
                12'd2020: logsin <= 24'd00691986;
                12'd2021: logsin <= 24'd00692674;
                12'd2022: logsin <= 24'd00693362;
                12'd2023: logsin <= 24'd00694050;
                12'd2024: logsin <= 24'd00694738;
                12'd2025: logsin <= 24'd00695427;
                12'd2026: logsin <= 24'd00696116;
                12'd2027: logsin <= 24'd00696806;
                12'd2028: logsin <= 24'd00697495;
                12'd2029: logsin <= 24'd00698185;
                12'd2030: logsin <= 24'd00698876;
                12'd2031: logsin <= 24'd00699566;
                12'd2032: logsin <= 24'd00700257;
                12'd2033: logsin <= 24'd00700949;
                12'd2034: logsin <= 24'd00701641;
                12'd2035: logsin <= 24'd00702332;
                12'd2036: logsin <= 24'd00703025;
                12'd2037: logsin <= 24'd00703717;
                12'd2038: logsin <= 24'd00704410;
                12'd2039: logsin <= 24'd00705104;
                12'd2040: logsin <= 24'd00705797;
                12'd2041: logsin <= 24'd00706491;
                12'd2042: logsin <= 24'd00707185;
                12'd2043: logsin <= 24'd00707880;
                12'd2044: logsin <= 24'd00708575;
                12'd2045: logsin <= 24'd00709270;
                12'd2046: logsin <= 24'd00709966;
                12'd2047: logsin <= 24'd00710662;
                12'd2048: logsin <= 24'd00711358;
                12'd2049: logsin <= 24'd00712054;
                12'd2050: logsin <= 24'd00712751;
                12'd2051: logsin <= 24'd00713448;
                12'd2052: logsin <= 24'd00714146;
                12'd2053: logsin <= 24'd00714843;
                12'd2054: logsin <= 24'd00715541;
                12'd2055: logsin <= 24'd00716240;
                12'd2056: logsin <= 24'd00716939;
                12'd2057: logsin <= 24'd00717638;
                12'd2058: logsin <= 24'd00718337;
                12'd2059: logsin <= 24'd00719037;
                12'd2060: logsin <= 24'd00719737;
                12'd2061: logsin <= 24'd00720437;
                12'd2062: logsin <= 24'd00721138;
                12'd2063: logsin <= 24'd00721839;
                12'd2064: logsin <= 24'd00722540;
                12'd2065: logsin <= 24'd00723242;
                12'd2066: logsin <= 24'd00723943;
                12'd2067: logsin <= 24'd00724646;
                12'd2068: logsin <= 24'd00725348;
                12'd2069: logsin <= 24'd00726051;
                12'd2070: logsin <= 24'd00726754;
                12'd2071: logsin <= 24'd00727458;
                12'd2072: logsin <= 24'd00728162;
                12'd2073: logsin <= 24'd00728866;
                12'd2074: logsin <= 24'd00729570;
                12'd2075: logsin <= 24'd00730275;
                12'd2076: logsin <= 24'd00730980;
                12'd2077: logsin <= 24'd00731685;
                12'd2078: logsin <= 24'd00732391;
                12'd2079: logsin <= 24'd00733097;
                12'd2080: logsin <= 24'd00733804;
                12'd2081: logsin <= 24'd00734510;
                12'd2082: logsin <= 24'd00735217;
                12'd2083: logsin <= 24'd00735925;
                12'd2084: logsin <= 24'd00736632;
                12'd2085: logsin <= 24'd00737340;
                12'd2086: logsin <= 24'd00738048;
                12'd2087: logsin <= 24'd00738757;
                12'd2088: logsin <= 24'd00739466;
                12'd2089: logsin <= 24'd00740175;
                12'd2090: logsin <= 24'd00740885;
                12'd2091: logsin <= 24'd00741594;
                12'd2092: logsin <= 24'd00742305;
                12'd2093: logsin <= 24'd00743015;
                12'd2094: logsin <= 24'd00743726;
                12'd2095: logsin <= 24'd00744437;
                12'd2096: logsin <= 24'd00745148;
                12'd2097: logsin <= 24'd00745860;
                12'd2098: logsin <= 24'd00746572;
                12'd2099: logsin <= 24'd00747284;
                12'd2100: logsin <= 24'd00747997;
                12'd2101: logsin <= 24'd00748710;
                12'd2102: logsin <= 24'd00749423;
                12'd2103: logsin <= 24'd00750137;
                12'd2104: logsin <= 24'd00750851;
                12'd2105: logsin <= 24'd00751565;
                12'd2106: logsin <= 24'd00752280;
                12'd2107: logsin <= 24'd00752995;
                12'd2108: logsin <= 24'd00753710;
                12'd2109: logsin <= 24'd00754425;
                12'd2110: logsin <= 24'd00755141;
                12'd2111: logsin <= 24'd00755857;
                12'd2112: logsin <= 24'd00756574;
                12'd2113: logsin <= 24'd00757290;
                12'd2114: logsin <= 24'd00758007;
                12'd2115: logsin <= 24'd00758725;
                12'd2116: logsin <= 24'd00759442;
                12'd2117: logsin <= 24'd00760160;
                12'd2118: logsin <= 24'd00760879;
                12'd2119: logsin <= 24'd00761597;
                12'd2120: logsin <= 24'd00762316;
                12'd2121: logsin <= 24'd00763035;
                12'd2122: logsin <= 24'd00763755;
                12'd2123: logsin <= 24'd00764475;
                12'd2124: logsin <= 24'd00765195;
                12'd2125: logsin <= 24'd00765915;
                12'd2126: logsin <= 24'd00766636;
                12'd2127: logsin <= 24'd00767357;
                12'd2128: logsin <= 24'd00768079;
                12'd2129: logsin <= 24'd00768800;
                12'd2130: logsin <= 24'd00769522;
                12'd2131: logsin <= 24'd00770245;
                12'd2132: logsin <= 24'd00770967;
                12'd2133: logsin <= 24'd00771690;
                12'd2134: logsin <= 24'd00772414;
                12'd2135: logsin <= 24'd00773137;
                12'd2136: logsin <= 24'd00773861;
                12'd2137: logsin <= 24'd00774585;
                12'd2138: logsin <= 24'd00775310;
                12'd2139: logsin <= 24'd00776035;
                12'd2140: logsin <= 24'd00776760;
                12'd2141: logsin <= 24'd00777485;
                12'd2142: logsin <= 24'd00778211;
                12'd2143: logsin <= 24'd00778937;
                12'd2144: logsin <= 24'd00779663;
                12'd2145: logsin <= 24'd00780390;
                12'd2146: logsin <= 24'd00781117;
                12'd2147: logsin <= 24'd00781844;
                12'd2148: logsin <= 24'd00782572;
                12'd2149: logsin <= 24'd00783300;
                12'd2150: logsin <= 24'd00784028;
                12'd2151: logsin <= 24'd00784756;
                12'd2152: logsin <= 24'd00785485;
                12'd2153: logsin <= 24'd00786214;
                12'd2154: logsin <= 24'd00786944;
                12'd2155: logsin <= 24'd00787673;
                12'd2156: logsin <= 24'd00788403;
                12'd2157: logsin <= 24'd00789134;
                12'd2158: logsin <= 24'd00789864;
                12'd2159: logsin <= 24'd00790595;
                12'd2160: logsin <= 24'd00791326;
                12'd2161: logsin <= 24'd00792058;
                12'd2162: logsin <= 24'd00792790;
                12'd2163: logsin <= 24'd00793522;
                12'd2164: logsin <= 24'd00794255;
                12'd2165: logsin <= 24'd00794987;
                12'd2166: logsin <= 24'd00795720;
                12'd2167: logsin <= 24'd00796454;
                12'd2168: logsin <= 24'd00797187;
                12'd2169: logsin <= 24'd00797921;
                12'd2170: logsin <= 24'd00798656;
                12'd2171: logsin <= 24'd00799390;
                12'd2172: logsin <= 24'd00800125;
                12'd2173: logsin <= 24'd00800860;
                12'd2174: logsin <= 24'd00801596;
                12'd2175: logsin <= 24'd00802332;
                12'd2176: logsin <= 24'd00803068;
                12'd2177: logsin <= 24'd00803804;
                12'd2178: logsin <= 24'd00804541;
                12'd2179: logsin <= 24'd00805278;
                12'd2180: logsin <= 24'd00806015;
                12'd2181: logsin <= 24'd00806753;
                12'd2182: logsin <= 24'd00807491;
                12'd2183: logsin <= 24'd00808229;
                12'd2184: logsin <= 24'd00808968;
                12'd2185: logsin <= 24'd00809706;
                12'd2186: logsin <= 24'd00810446;
                12'd2187: logsin <= 24'd00811185;
                12'd2188: logsin <= 24'd00811925;
                12'd2189: logsin <= 24'd00812665;
                12'd2190: logsin <= 24'd00813405;
                12'd2191: logsin <= 24'd00814146;
                12'd2192: logsin <= 24'd00814887;
                12'd2193: logsin <= 24'd00815628;
                12'd2194: logsin <= 24'd00816369;
                12'd2195: logsin <= 24'd00817111;
                12'd2196: logsin <= 24'd00817853;
                12'd2197: logsin <= 24'd00818596;
                12'd2198: logsin <= 24'd00819338;
                12'd2199: logsin <= 24'd00820081;
                12'd2200: logsin <= 24'd00820825;
                12'd2201: logsin <= 24'd00821568;
                12'd2202: logsin <= 24'd00822312;
                12'd2203: logsin <= 24'd00823057;
                12'd2204: logsin <= 24'd00823801;
                12'd2205: logsin <= 24'd00824546;
                12'd2206: logsin <= 24'd00825291;
                12'd2207: logsin <= 24'd00826036;
                12'd2208: logsin <= 24'd00826782;
                12'd2209: logsin <= 24'd00827528;
                12'd2210: logsin <= 24'd00828274;
                12'd2211: logsin <= 24'd00829021;
                12'd2212: logsin <= 24'd00829768;
                12'd2213: logsin <= 24'd00830515;
                12'd2214: logsin <= 24'd00831263;
                12'd2215: logsin <= 24'd00832010;
                12'd2216: logsin <= 24'd00832758;
                12'd2217: logsin <= 24'd00833507;
                12'd2218: logsin <= 24'd00834255;
                12'd2219: logsin <= 24'd00835004;
                12'd2220: logsin <= 24'd00835754;
                12'd2221: logsin <= 24'd00836503;
                12'd2222: logsin <= 24'd00837253;
                12'd2223: logsin <= 24'd00838003;
                12'd2224: logsin <= 24'd00838754;
                12'd2225: logsin <= 24'd00839504;
                12'd2226: logsin <= 24'd00840255;
                12'd2227: logsin <= 24'd00841007;
                12'd2228: logsin <= 24'd00841758;
                12'd2229: logsin <= 24'd00842510;
                12'd2230: logsin <= 24'd00843262;
                12'd2231: logsin <= 24'd00844015;
                12'd2232: logsin <= 24'd00844768;
                12'd2233: logsin <= 24'd00845521;
                12'd2234: logsin <= 24'd00846274;
                12'd2235: logsin <= 24'd00847028;
                12'd2236: logsin <= 24'd00847782;
                12'd2237: logsin <= 24'd00848536;
                12'd2238: logsin <= 24'd00849290;
                12'd2239: logsin <= 24'd00850045;
                12'd2240: logsin <= 24'd00850800;
                12'd2241: logsin <= 24'd00851556;
                12'd2242: logsin <= 24'd00852312;
                12'd2243: logsin <= 24'd00853067;
                12'd2244: logsin <= 24'd00853824;
                12'd2245: logsin <= 24'd00854580;
                12'd2246: logsin <= 24'd00855337;
                12'd2247: logsin <= 24'd00856094;
                12'd2248: logsin <= 24'd00856852;
                12'd2249: logsin <= 24'd00857610;
                12'd2250: logsin <= 24'd00858368;
                12'd2251: logsin <= 24'd00859126;
                12'd2252: logsin <= 24'd00859884;
                12'd2253: logsin <= 24'd00860643;
                12'd2254: logsin <= 24'd00861402;
                12'd2255: logsin <= 24'd00862162;
                12'd2256: logsin <= 24'd00862922;
                12'd2257: logsin <= 24'd00863682;
                12'd2258: logsin <= 24'd00864442;
                12'd2259: logsin <= 24'd00865203;
                12'd2260: logsin <= 24'd00865964;
                12'd2261: logsin <= 24'd00866725;
                12'd2262: logsin <= 24'd00867486;
                12'd2263: logsin <= 24'd00868248;
                12'd2264: logsin <= 24'd00869010;
                12'd2265: logsin <= 24'd00869772;
                12'd2266: logsin <= 24'd00870535;
                12'd2267: logsin <= 24'd00871298;
                12'd2268: logsin <= 24'd00872061;
                12'd2269: logsin <= 24'd00872824;
                12'd2270: logsin <= 24'd00873588;
                12'd2271: logsin <= 24'd00874352;
                12'd2272: logsin <= 24'd00875117;
                12'd2273: logsin <= 24'd00875881;
                12'd2274: logsin <= 24'd00876646;
                12'd2275: logsin <= 24'd00877411;
                12'd2276: logsin <= 24'd00878177;
                12'd2277: logsin <= 24'd00878942;
                12'd2278: logsin <= 24'd00879708;
                12'd2279: logsin <= 24'd00880475;
                12'd2280: logsin <= 24'd00881241;
                12'd2281: logsin <= 24'd00882008;
                12'd2282: logsin <= 24'd00882775;
                12'd2283: logsin <= 24'd00883543;
                12'd2284: logsin <= 24'd00884311;
                12'd2285: logsin <= 24'd00885079;
                12'd2286: logsin <= 24'd00885847;
                12'd2287: logsin <= 24'd00886615;
                12'd2288: logsin <= 24'd00887384;
                12'd2289: logsin <= 24'd00888153;
                12'd2290: logsin <= 24'd00888923;
                12'd2291: logsin <= 24'd00889692;
                12'd2292: logsin <= 24'd00890462;
                12'd2293: logsin <= 24'd00891233;
                12'd2294: logsin <= 24'd00892003;
                12'd2295: logsin <= 24'd00892774;
                12'd2296: logsin <= 24'd00893545;
                12'd2297: logsin <= 24'd00894317;
                12'd2298: logsin <= 24'd00895088;
                12'd2299: logsin <= 24'd00895860;
                12'd2300: logsin <= 24'd00896632;
                12'd2301: logsin <= 24'd00897405;
                12'd2302: logsin <= 24'd00898178;
                12'd2303: logsin <= 24'd00898951;
                12'd2304: logsin <= 24'd00899724;
                12'd2305: logsin <= 24'd00900497;
                12'd2306: logsin <= 24'd00901271;
                12'd2307: logsin <= 24'd00902045;
                12'd2308: logsin <= 24'd00902820;
                12'd2309: logsin <= 24'd00903595;
                12'd2310: logsin <= 24'd00904370;
                12'd2311: logsin <= 24'd00905145;
                12'd2312: logsin <= 24'd00905920;
                12'd2313: logsin <= 24'd00906696;
                12'd2314: logsin <= 24'd00907472;
                12'd2315: logsin <= 24'd00908249;
                12'd2316: logsin <= 24'd00909025;
                12'd2317: logsin <= 24'd00909802;
                12'd2318: logsin <= 24'd00910579;
                12'd2319: logsin <= 24'd00911357;
                12'd2320: logsin <= 24'd00912134;
                12'd2321: logsin <= 24'd00912912;
                12'd2322: logsin <= 24'd00913691;
                12'd2323: logsin <= 24'd00914469;
                12'd2324: logsin <= 24'd00915248;
                12'd2325: logsin <= 24'd00916027;
                12'd2326: logsin <= 24'd00916806;
                12'd2327: logsin <= 24'd00917586;
                12'd2328: logsin <= 24'd00918366;
                12'd2329: logsin <= 24'd00919146;
                12'd2330: logsin <= 24'd00919927;
                12'd2331: logsin <= 24'd00920707;
                12'd2332: logsin <= 24'd00921488;
                12'd2333: logsin <= 24'd00922270;
                12'd2334: logsin <= 24'd00923051;
                12'd2335: logsin <= 24'd00923833;
                12'd2336: logsin <= 24'd00924615;
                12'd2337: logsin <= 24'd00925397;
                12'd2338: logsin <= 24'd00926180;
                12'd2339: logsin <= 24'd00926963;
                12'd2340: logsin <= 24'd00927746;
                12'd2341: logsin <= 24'd00928529;
                12'd2342: logsin <= 24'd00929313;
                12'd2343: logsin <= 24'd00930097;
                12'd2344: logsin <= 24'd00930881;
                12'd2345: logsin <= 24'd00931666;
                12'd2346: logsin <= 24'd00932450;
                12'd2347: logsin <= 24'd00933235;
                12'd2348: logsin <= 24'd00934021;
                12'd2349: logsin <= 24'd00934806;
                12'd2350: logsin <= 24'd00935592;
                12'd2351: logsin <= 24'd00936378;
                12'd2352: logsin <= 24'd00937165;
                12'd2353: logsin <= 24'd00937951;
                12'd2354: logsin <= 24'd00938738;
                12'd2355: logsin <= 24'd00939525;
                12'd2356: logsin <= 24'd00940313;
                12'd2357: logsin <= 24'd00941100;
                12'd2358: logsin <= 24'd00941888;
                12'd2359: logsin <= 24'd00942676;
                12'd2360: logsin <= 24'd00943465;
                12'd2361: logsin <= 24'd00944254;
                12'd2362: logsin <= 24'd00945043;
                12'd2363: logsin <= 24'd00945832;
                12'd2364: logsin <= 24'd00946621;
                12'd2365: logsin <= 24'd00947411;
                12'd2366: logsin <= 24'd00948201;
                12'd2367: logsin <= 24'd00948991;
                12'd2368: logsin <= 24'd00949782;
                12'd2369: logsin <= 24'd00950573;
                12'd2370: logsin <= 24'd00951364;
                12'd2371: logsin <= 24'd00952155;
                12'd2372: logsin <= 24'd00952947;
                12'd2373: logsin <= 24'd00953739;
                12'd2374: logsin <= 24'd00954531;
                12'd2375: logsin <= 24'd00955323;
                12'd2376: logsin <= 24'd00956116;
                12'd2377: logsin <= 24'd00956909;
                12'd2378: logsin <= 24'd00957702;
                12'd2379: logsin <= 24'd00958495;
                12'd2380: logsin <= 24'd00959289;
                12'd2381: logsin <= 24'd00960083;
                12'd2382: logsin <= 24'd00960877;
                12'd2383: logsin <= 24'd00961672;
                12'd2384: logsin <= 24'd00962466;
                12'd2385: logsin <= 24'd00963261;
                12'd2386: logsin <= 24'd00964056;
                12'd2387: logsin <= 24'd00964852;
                12'd2388: logsin <= 24'd00965648;
                12'd2389: logsin <= 24'd00966444;
                12'd2390: logsin <= 24'd00967240;
                12'd2391: logsin <= 24'd00968036;
                12'd2392: logsin <= 24'd00968833;
                12'd2393: logsin <= 24'd00969630;
                12'd2394: logsin <= 24'd00970427;
                12'd2395: logsin <= 24'd00971225;
                12'd2396: logsin <= 24'd00972023;
                12'd2397: logsin <= 24'd00972821;
                12'd2398: logsin <= 24'd00973619;
                12'd2399: logsin <= 24'd00974418;
                12'd2400: logsin <= 24'd00975216;
                12'd2401: logsin <= 24'd00976015;
                12'd2402: logsin <= 24'd00976815;
                12'd2403: logsin <= 24'd00977614;
                12'd2404: logsin <= 24'd00978414;
                12'd2405: logsin <= 24'd00979214;
                12'd2406: logsin <= 24'd00980014;
                12'd2407: logsin <= 24'd00980815;
                12'd2408: logsin <= 24'd00981616;
                12'd2409: logsin <= 24'd00982417;
                12'd2410: logsin <= 24'd00983218;
                12'd2411: logsin <= 24'd00984019;
                12'd2412: logsin <= 24'd00984821;
                12'd2413: logsin <= 24'd00985623;
                12'd2414: logsin <= 24'd00986426;
                12'd2415: logsin <= 24'd00987228;
                12'd2416: logsin <= 24'd00988031;
                12'd2417: logsin <= 24'd00988834;
                12'd2418: logsin <= 24'd00989637;
                12'd2419: logsin <= 24'd00990441;
                12'd2420: logsin <= 24'd00991244;
                12'd2421: logsin <= 24'd00992048;
                12'd2422: logsin <= 24'd00992853;
                12'd2423: logsin <= 24'd00993657;
                12'd2424: logsin <= 24'd00994462;
                12'd2425: logsin <= 24'd00995267;
                12'd2426: logsin <= 24'd00996072;
                12'd2427: logsin <= 24'd00996878;
                12'd2428: logsin <= 24'd00997683;
                12'd2429: logsin <= 24'd00998489;
                12'd2430: logsin <= 24'd00999296;
                12'd2431: logsin <= 24'd01000102;
                12'd2432: logsin <= 24'd01000909;
                12'd2433: logsin <= 24'd01001716;
                12'd2434: logsin <= 24'd01002523;
                12'd2435: logsin <= 24'd01003330;
                12'd2436: logsin <= 24'd01004138;
                12'd2437: logsin <= 24'd01004946;
                12'd2438: logsin <= 24'd01005754;
                12'd2439: logsin <= 24'd01006562;
                12'd2440: logsin <= 24'd01007371;
                12'd2441: logsin <= 24'd01008180;
                12'd2442: logsin <= 24'd01008989;
                12'd2443: logsin <= 24'd01009798;
                12'd2444: logsin <= 24'd01010608;
                12'd2445: logsin <= 24'd01011418;
                12'd2446: logsin <= 24'd01012228;
                12'd2447: logsin <= 24'd01013038;
                12'd2448: logsin <= 24'd01013849;
                12'd2449: logsin <= 24'd01014659;
                12'd2450: logsin <= 24'd01015470;
                12'd2451: logsin <= 24'd01016282;
                12'd2452: logsin <= 24'd01017093;
                12'd2453: logsin <= 24'd01017905;
                12'd2454: logsin <= 24'd01018717;
                12'd2455: logsin <= 24'd01019529;
                12'd2456: logsin <= 24'd01020341;
                12'd2457: logsin <= 24'd01021154;
                12'd2458: logsin <= 24'd01021967;
                12'd2459: logsin <= 24'd01022780;
                12'd2460: logsin <= 24'd01023593;
                12'd2461: logsin <= 24'd01024407;
                12'd2462: logsin <= 24'd01025221;
                12'd2463: logsin <= 24'd01026035;
                12'd2464: logsin <= 24'd01026849;
                12'd2465: logsin <= 24'd01027664;
                12'd2466: logsin <= 24'd01028478;
                12'd2467: logsin <= 24'd01029293;
                12'd2468: logsin <= 24'd01030109;
                12'd2469: logsin <= 24'd01030924;
                12'd2470: logsin <= 24'd01031740;
                12'd2471: logsin <= 24'd01032556;
                12'd2472: logsin <= 24'd01033372;
                12'd2473: logsin <= 24'd01034188;
                12'd2474: logsin <= 24'd01035005;
                12'd2475: logsin <= 24'd01035822;
                12'd2476: logsin <= 24'd01036639;
                12'd2477: logsin <= 24'd01037456;
                12'd2478: logsin <= 24'd01038273;
                12'd2479: logsin <= 24'd01039091;
                12'd2480: logsin <= 24'd01039909;
                12'd2481: logsin <= 24'd01040727;
                12'd2482: logsin <= 24'd01041546;
                12'd2483: logsin <= 24'd01042364;
                12'd2484: logsin <= 24'd01043183;
                12'd2485: logsin <= 24'd01044002;
                12'd2486: logsin <= 24'd01044822;
                12'd2487: logsin <= 24'd01045641;
                12'd2488: logsin <= 24'd01046461;
                12'd2489: logsin <= 24'd01047281;
                12'd2490: logsin <= 24'd01048101;
                12'd2491: logsin <= 24'd01048922;
                12'd2492: logsin <= 24'd01049742;
                12'd2493: logsin <= 24'd01050563;
                12'd2494: logsin <= 24'd01051384;
                12'd2495: logsin <= 24'd01052205;
                12'd2496: logsin <= 24'd01053027;
                12'd2497: logsin <= 24'd01053849;
                12'd2498: logsin <= 24'd01054671;
                12'd2499: logsin <= 24'd01055493;
                12'd2500: logsin <= 24'd01056315;
                12'd2501: logsin <= 24'd01057138;
                12'd2502: logsin <= 24'd01057961;
                12'd2503: logsin <= 24'd01058784;
                12'd2504: logsin <= 24'd01059607;
                12'd2505: logsin <= 24'd01060431;
                12'd2506: logsin <= 24'd01061254;
                12'd2507: logsin <= 24'd01062078;
                12'd2508: logsin <= 24'd01062903;
                12'd2509: logsin <= 24'd01063727;
                12'd2510: logsin <= 24'd01064551;
                12'd2511: logsin <= 24'd01065376;
                12'd2512: logsin <= 24'd01066201;
                12'd2513: logsin <= 24'd01067027;
                12'd2514: logsin <= 24'd01067852;
                12'd2515: logsin <= 24'd01068678;
                12'd2516: logsin <= 24'd01069504;
                12'd2517: logsin <= 24'd01070330;
                12'd2518: logsin <= 24'd01071156;
                12'd2519: logsin <= 24'd01071982;
                12'd2520: logsin <= 24'd01072809;
                12'd2521: logsin <= 24'd01073636;
                12'd2522: logsin <= 24'd01074463;
                12'd2523: logsin <= 24'd01075291;
                12'd2524: logsin <= 24'd01076118;
                12'd2525: logsin <= 24'd01076946;
                12'd2526: logsin <= 24'd01077774;
                12'd2527: logsin <= 24'd01078602;
                12'd2528: logsin <= 24'd01079431;
                12'd2529: logsin <= 24'd01080259;
                12'd2530: logsin <= 24'd01081088;
                12'd2531: logsin <= 24'd01081917;
                12'd2532: logsin <= 24'd01082746;
                12'd2533: logsin <= 24'd01083576;
                12'd2534: logsin <= 24'd01084405;
                12'd2535: logsin <= 24'd01085235;
                12'd2536: logsin <= 24'd01086065;
                12'd2537: logsin <= 24'd01086895;
                12'd2538: logsin <= 24'd01087726;
                12'd2539: logsin <= 24'd01088557;
                12'd2540: logsin <= 24'd01089388;
                12'd2541: logsin <= 24'd01090219;
                12'd2542: logsin <= 24'd01091050;
                12'd2543: logsin <= 24'd01091881;
                12'd2544: logsin <= 24'd01092713;
                12'd2545: logsin <= 24'd01093545;
                12'd2546: logsin <= 24'd01094377;
                12'd2547: logsin <= 24'd01095209;
                12'd2548: logsin <= 24'd01096042;
                12'd2549: logsin <= 24'd01096875;
                12'd2550: logsin <= 24'd01097707;
                12'd2551: logsin <= 24'd01098541;
                12'd2552: logsin <= 24'd01099374;
                12'd2553: logsin <= 24'd01100207;
                12'd2554: logsin <= 24'd01101041;
                12'd2555: logsin <= 24'd01101875;
                12'd2556: logsin <= 24'd01102709;
                12'd2557: logsin <= 24'd01103543;
                12'd2558: logsin <= 24'd01104378;
                12'd2559: logsin <= 24'd01105212;
                12'd2560: logsin <= 24'd01106047;
                12'd2561: logsin <= 24'd01106882;
                12'd2562: logsin <= 24'd01107718;
                12'd2563: logsin <= 24'd01108553;
                12'd2564: logsin <= 24'd01109389;
                12'd2565: logsin <= 24'd01110225;
                12'd2566: logsin <= 24'd01111061;
                12'd2567: logsin <= 24'd01111897;
                12'd2568: logsin <= 24'd01112733;
                12'd2569: logsin <= 24'd01113570;
                12'd2570: logsin <= 24'd01114407;
                12'd2571: logsin <= 24'd01115244;
                12'd2572: logsin <= 24'd01116081;
                12'd2573: logsin <= 24'd01116918;
                12'd2574: logsin <= 24'd01117756;
                12'd2575: logsin <= 24'd01118594;
                12'd2576: logsin <= 24'd01119432;
                12'd2577: logsin <= 24'd01120270;
                12'd2578: logsin <= 24'd01121108;
                12'd2579: logsin <= 24'd01121947;
                12'd2580: logsin <= 24'd01122785;
                12'd2581: logsin <= 24'd01123624;
                12'd2582: logsin <= 24'd01124463;
                12'd2583: logsin <= 24'd01125302;
                12'd2584: logsin <= 24'd01126142;
                12'd2585: logsin <= 24'd01126981;
                12'd2586: logsin <= 24'd01127821;
                12'd2587: logsin <= 24'd01128661;
                12'd2588: logsin <= 24'd01129501;
                12'd2589: logsin <= 24'd01130342;
                12'd2590: logsin <= 24'd01131182;
                12'd2591: logsin <= 24'd01132023;
                12'd2592: logsin <= 24'd01132864;
                12'd2593: logsin <= 24'd01133705;
                12'd2594: logsin <= 24'd01134546;
                12'd2595: logsin <= 24'd01135388;
                12'd2596: logsin <= 24'd01136229;
                12'd2597: logsin <= 24'd01137071;
                12'd2598: logsin <= 24'd01137913;
                12'd2599: logsin <= 24'd01138755;
                12'd2600: logsin <= 24'd01139598;
                12'd2601: logsin <= 24'd01140440;
                12'd2602: logsin <= 24'd01141283;
                12'd2603: logsin <= 24'd01142126;
                12'd2604: logsin <= 24'd01142969;
                12'd2605: logsin <= 24'd01143812;
                12'd2606: logsin <= 24'd01144656;
                12'd2607: logsin <= 24'd01145499;
                12'd2608: logsin <= 24'd01146343;
                12'd2609: logsin <= 24'd01147187;
                12'd2610: logsin <= 24'd01148031;
                12'd2611: logsin <= 24'd01148875;
                12'd2612: logsin <= 24'd01149720;
                12'd2613: logsin <= 24'd01150564;
                12'd2614: logsin <= 24'd01151409;
                12'd2615: logsin <= 24'd01152254;
                12'd2616: logsin <= 24'd01153099;
                12'd2617: logsin <= 24'd01153944;
                12'd2618: logsin <= 24'd01154790;
                12'd2619: logsin <= 24'd01155636;
                12'd2620: logsin <= 24'd01156481;
                12'd2621: logsin <= 24'd01157327;
                12'd2622: logsin <= 24'd01158174;
                12'd2623: logsin <= 24'd01159020;
                12'd2624: logsin <= 24'd01159866;
                12'd2625: logsin <= 24'd01160713;
                12'd2626: logsin <= 24'd01161560;
                12'd2627: logsin <= 24'd01162407;
                12'd2628: logsin <= 24'd01163254;
                12'd2629: logsin <= 24'd01164101;
                12'd2630: logsin <= 24'd01164949;
                12'd2631: logsin <= 24'd01165796;
                12'd2632: logsin <= 24'd01166644;
                12'd2633: logsin <= 24'd01167492;
                12'd2634: logsin <= 24'd01168340;
                12'd2635: logsin <= 24'd01169188;
                12'd2636: logsin <= 24'd01170037;
                12'd2637: logsin <= 24'd01170886;
                12'd2638: logsin <= 24'd01171734;
                12'd2639: logsin <= 24'd01172583;
                12'd2640: logsin <= 24'd01173432;
                12'd2641: logsin <= 24'd01174282;
                12'd2642: logsin <= 24'd01175131;
                12'd2643: logsin <= 24'd01175980;
                12'd2644: logsin <= 24'd01176830;
                12'd2645: logsin <= 24'd01177680;
                12'd2646: logsin <= 24'd01178530;
                12'd2647: logsin <= 24'd01179380;
                12'd2648: logsin <= 24'd01180231;
                12'd2649: logsin <= 24'd01181081;
                12'd2650: logsin <= 24'd01181932;
                12'd2651: logsin <= 24'd01182783;
                12'd2652: logsin <= 24'd01183634;
                12'd2653: logsin <= 24'd01184485;
                12'd2654: logsin <= 24'd01185336;
                12'd2655: logsin <= 24'd01186187;
                12'd2656: logsin <= 24'd01187039;
                12'd2657: logsin <= 24'd01187891;
                12'd2658: logsin <= 24'd01188742;
                12'd2659: logsin <= 24'd01189594;
                12'd2660: logsin <= 24'd01190447;
                12'd2661: logsin <= 24'd01191299;
                12'd2662: logsin <= 24'd01192151;
                12'd2663: logsin <= 24'd01193004;
                12'd2664: logsin <= 24'd01193857;
                12'd2665: logsin <= 24'd01194710;
                12'd2666: logsin <= 24'd01195563;
                12'd2667: logsin <= 24'd01196416;
                12'd2668: logsin <= 24'd01197269;
                12'd2669: logsin <= 24'd01198123;
                12'd2670: logsin <= 24'd01198976;
                12'd2671: logsin <= 24'd01199830;
                12'd2672: logsin <= 24'd01200684;
                12'd2673: logsin <= 24'd01201538;
                12'd2674: logsin <= 24'd01202392;
                12'd2675: logsin <= 24'd01203246;
                12'd2676: logsin <= 24'd01204101;
                12'd2677: logsin <= 24'd01204956;
                12'd2678: logsin <= 24'd01205810;
                12'd2679: logsin <= 24'd01206665;
                12'd2680: logsin <= 24'd01207520;
                12'd2681: logsin <= 24'd01208375;
                12'd2682: logsin <= 24'd01209231;
                12'd2683: logsin <= 24'd01210086;
                12'd2684: logsin <= 24'd01210942;
                12'd2685: logsin <= 24'd01211797;
                12'd2686: logsin <= 24'd01212653;
                12'd2687: logsin <= 24'd01213509;
                12'd2688: logsin <= 24'd01214365;
                12'd2689: logsin <= 24'd01215221;
                12'd2690: logsin <= 24'd01216078;
                12'd2691: logsin <= 24'd01216934;
                12'd2692: logsin <= 24'd01217791;
                12'd2693: logsin <= 24'd01218648;
                12'd2694: logsin <= 24'd01219505;
                12'd2695: logsin <= 24'd01220362;
                12'd2696: logsin <= 24'd01221219;
                12'd2697: logsin <= 24'd01222076;
                12'd2698: logsin <= 24'd01222934;
                12'd2699: logsin <= 24'd01223791;
                12'd2700: logsin <= 24'd01224649;
                12'd2701: logsin <= 24'd01225507;
                12'd2702: logsin <= 24'd01226364;
                12'd2703: logsin <= 24'd01227223;
                12'd2704: logsin <= 24'd01228081;
                12'd2705: logsin <= 24'd01228939;
                12'd2706: logsin <= 24'd01229797;
                12'd2707: logsin <= 24'd01230656;
                12'd2708: logsin <= 24'd01231515;
                12'd2709: logsin <= 24'd01232373;
                12'd2710: logsin <= 24'd01233232;
                12'd2711: logsin <= 24'd01234091;
                12'd2712: logsin <= 24'd01234950;
                12'd2713: logsin <= 24'd01235810;
                12'd2714: logsin <= 24'd01236669;
                12'd2715: logsin <= 24'd01237529;
                12'd2716: logsin <= 24'd01238388;
                12'd2717: logsin <= 24'd01239248;
                12'd2718: logsin <= 24'd01240108;
                12'd2719: logsin <= 24'd01240968;
                12'd2720: logsin <= 24'd01241828;
                12'd2721: logsin <= 24'd01242688;
                12'd2722: logsin <= 24'd01243548;
                12'd2723: logsin <= 24'd01244409;
                12'd2724: logsin <= 24'd01245269;
                12'd2725: logsin <= 24'd01246130;
                12'd2726: logsin <= 24'd01246991;
                12'd2727: logsin <= 24'd01247852;
                12'd2728: logsin <= 24'd01248713;
                12'd2729: logsin <= 24'd01249574;
                12'd2730: logsin <= 24'd01250435;
                12'd2731: logsin <= 24'd01251296;
                12'd2732: logsin <= 24'd01252158;
                12'd2733: logsin <= 24'd01253019;
                12'd2734: logsin <= 24'd01253881;
                12'd2735: logsin <= 24'd01254743;
                12'd2736: logsin <= 24'd01255605;
                12'd2737: logsin <= 24'd01256467;
                12'd2738: logsin <= 24'd01257329;
                12'd2739: logsin <= 24'd01258191;
                12'd2740: logsin <= 24'd01259053;
                12'd2741: logsin <= 24'd01259916;
                12'd2742: logsin <= 24'd01260778;
                12'd2743: logsin <= 24'd01261641;
                12'd2744: logsin <= 24'd01262503;
                12'd2745: logsin <= 24'd01263366;
                12'd2746: logsin <= 24'd01264229;
                12'd2747: logsin <= 24'd01265092;
                12'd2748: logsin <= 24'd01265955;
                12'd2749: logsin <= 24'd01266818;
                12'd2750: logsin <= 24'd01267681;
                12'd2751: logsin <= 24'd01268545;
                12'd2752: logsin <= 24'd01269408;
                12'd2753: logsin <= 24'd01270272;
                12'd2754: logsin <= 24'd01271136;
                12'd2755: logsin <= 24'd01271999;
                12'd2756: logsin <= 24'd01272863;
                12'd2757: logsin <= 24'd01273727;
                12'd2758: logsin <= 24'd01274591;
                12'd2759: logsin <= 24'd01275455;
                12'd2760: logsin <= 24'd01276320;
                12'd2761: logsin <= 24'd01277184;
                12'd2762: logsin <= 24'd01278048;
                12'd2763: logsin <= 24'd01278913;
                12'd2764: logsin <= 24'd01279777;
                12'd2765: logsin <= 24'd01280642;
                12'd2766: logsin <= 24'd01281507;
                12'd2767: logsin <= 24'd01282372;
                12'd2768: logsin <= 24'd01283237;
                12'd2769: logsin <= 24'd01284102;
                12'd2770: logsin <= 24'd01284967;
                12'd2771: logsin <= 24'd01285832;
                12'd2772: logsin <= 24'd01286697;
                12'd2773: logsin <= 24'd01287562;
                12'd2774: logsin <= 24'd01288428;
                12'd2775: logsin <= 24'd01289293;
                12'd2776: logsin <= 24'd01290159;
                12'd2777: logsin <= 24'd01291025;
                12'd2778: logsin <= 24'd01291890;
                12'd2779: logsin <= 24'd01292756;
                12'd2780: logsin <= 24'd01293622;
                12'd2781: logsin <= 24'd01294488;
                12'd2782: logsin <= 24'd01295354;
                12'd2783: logsin <= 24'd01296220;
                12'd2784: logsin <= 24'd01297087;
                12'd2785: logsin <= 24'd01297953;
                12'd2786: logsin <= 24'd01298819;
                12'd2787: logsin <= 24'd01299686;
                12'd2788: logsin <= 24'd01300552;
                12'd2789: logsin <= 24'd01301419;
                12'd2790: logsin <= 24'd01302285;
                12'd2791: logsin <= 24'd01303152;
                12'd2792: logsin <= 24'd01304019;
                12'd2793: logsin <= 24'd01304886;
                12'd2794: logsin <= 24'd01305753;
                12'd2795: logsin <= 24'd01306620;
                12'd2796: logsin <= 24'd01307487;
                12'd2797: logsin <= 24'd01308354;
                12'd2798: logsin <= 24'd01309221;
                12'd2799: logsin <= 24'd01310088;
                12'd2800: logsin <= 24'd01310956;
                12'd2801: logsin <= 24'd01311823;
                12'd2802: logsin <= 24'd01312691;
                12'd2803: logsin <= 24'd01313558;
                12'd2804: logsin <= 24'd01314426;
                12'd2805: logsin <= 24'd01315293;
                12'd2806: logsin <= 24'd01316161;
                12'd2807: logsin <= 24'd01317029;
                12'd2808: logsin <= 24'd01317897;
                12'd2809: logsin <= 24'd01318765;
                12'd2810: logsin <= 24'd01319632;
                12'd2811: logsin <= 24'd01320500;
                12'd2812: logsin <= 24'd01321369;
                12'd2813: logsin <= 24'd01322237;
                12'd2814: logsin <= 24'd01323105;
                12'd2815: logsin <= 24'd01323973;
                12'd2816: logsin <= 24'd01324841;
                12'd2817: logsin <= 24'd01325710;
                12'd2818: logsin <= 24'd01326578;
                12'd2819: logsin <= 24'd01327446;
                12'd2820: logsin <= 24'd01328315;
                12'd2821: logsin <= 24'd01329184;
                12'd2822: logsin <= 24'd01330052;
                12'd2823: logsin <= 24'd01330921;
                12'd2824: logsin <= 24'd01331789;
                12'd2825: logsin <= 24'd01332658;
                12'd2826: logsin <= 24'd01333527;
                12'd2827: logsin <= 24'd01334396;
                12'd2828: logsin <= 24'd01335265;
                12'd2829: logsin <= 24'd01336134;
                12'd2830: logsin <= 24'd01337002;
                12'd2831: logsin <= 24'd01337871;
                12'd2832: logsin <= 24'd01338741;
                12'd2833: logsin <= 24'd01339610;
                12'd2834: logsin <= 24'd01340479;
                12'd2835: logsin <= 24'd01341348;
                12'd2836: logsin <= 24'd01342217;
                12'd2837: logsin <= 24'd01343086;
                12'd2838: logsin <= 24'd01343956;
                12'd2839: logsin <= 24'd01344825;
                12'd2840: logsin <= 24'd01345694;
                12'd2841: logsin <= 24'd01346564;
                12'd2842: logsin <= 24'd01347433;
                12'd2843: logsin <= 24'd01348303;
                12'd2844: logsin <= 24'd01349172;
                12'd2845: logsin <= 24'd01350042;
                12'd2846: logsin <= 24'd01350911;
                12'd2847: logsin <= 24'd01351781;
                12'd2848: logsin <= 24'd01352650;
                12'd2849: logsin <= 24'd01353520;
                12'd2850: logsin <= 24'd01354390;
                12'd2851: logsin <= 24'd01355259;
                12'd2852: logsin <= 24'd01356129;
                12'd2853: logsin <= 24'd01356999;
                12'd2854: logsin <= 24'd01357869;
                12'd2855: logsin <= 24'd01358738;
                12'd2856: logsin <= 24'd01359608;
                12'd2857: logsin <= 24'd01360478;
                12'd2858: logsin <= 24'd01361348;
                12'd2859: logsin <= 24'd01362218;
                12'd2860: logsin <= 24'd01363088;
                12'd2861: logsin <= 24'd01363958;
                12'd2862: logsin <= 24'd01364828;
                12'd2863: logsin <= 24'd01365698;
                12'd2864: logsin <= 24'd01366568;
                12'd2865: logsin <= 24'd01367438;
                12'd2866: logsin <= 24'd01368308;
                12'd2867: logsin <= 24'd01369178;
                12'd2868: logsin <= 24'd01370048;
                12'd2869: logsin <= 24'd01370918;
                12'd2870: logsin <= 24'd01371788;
                12'd2871: logsin <= 24'd01372658;
                12'd2872: logsin <= 24'd01373528;
                12'd2873: logsin <= 24'd01374399;
                12'd2874: logsin <= 24'd01375269;
                12'd2875: logsin <= 24'd01376139;
                12'd2876: logsin <= 24'd01377009;
                12'd2877: logsin <= 24'd01377879;
                12'd2878: logsin <= 24'd01378749;
                12'd2879: logsin <= 24'd01379620;
                12'd2880: logsin <= 24'd01380490;
                12'd2881: logsin <= 24'd01381360;
                12'd2882: logsin <= 24'd01382230;
                12'd2883: logsin <= 24'd01383100;
                12'd2884: logsin <= 24'd01383971;
                12'd2885: logsin <= 24'd01384841;
                12'd2886: logsin <= 24'd01385711;
                12'd2887: logsin <= 24'd01386581;
                12'd2888: logsin <= 24'd01387451;
                12'd2889: logsin <= 24'd01388322;
                12'd2890: logsin <= 24'd01389192;
                12'd2891: logsin <= 24'd01390062;
                12'd2892: logsin <= 24'd01390932;
                12'd2893: logsin <= 24'd01391802;
                12'd2894: logsin <= 24'd01392673;
                12'd2895: logsin <= 24'd01393543;
                12'd2896: logsin <= 24'd01394413;
                12'd2897: logsin <= 24'd01395283;
                12'd2898: logsin <= 24'd01396153;
                12'd2899: logsin <= 24'd01397023;
                12'd2900: logsin <= 24'd01397894;
                12'd2901: logsin <= 24'd01398764;
                12'd2902: logsin <= 24'd01399634;
                12'd2903: logsin <= 24'd01400504;
                12'd2904: logsin <= 24'd01401374;
                12'd2905: logsin <= 24'd01402244;
                12'd2906: logsin <= 24'd01403114;
                12'd2907: logsin <= 24'd01403984;
                12'd2908: logsin <= 24'd01404854;
                12'd2909: logsin <= 24'd01405724;
                12'd2910: logsin <= 24'd01406594;
                12'd2911: logsin <= 24'd01407464;
                12'd2912: logsin <= 24'd01408334;
                12'd2913: logsin <= 24'd01409204;
                12'd2914: logsin <= 24'd01410074;
                12'd2915: logsin <= 24'd01410944;
                12'd2916: logsin <= 24'd01411814;
                12'd2917: logsin <= 24'd01412684;
                12'd2918: logsin <= 24'd01413554;
                12'd2919: logsin <= 24'd01414423;
                12'd2920: logsin <= 24'd01415293;
                12'd2921: logsin <= 24'd01416163;
                12'd2922: logsin <= 24'd01417033;
                12'd2923: logsin <= 24'd01417902;
                12'd2924: logsin <= 24'd01418772;
                12'd2925: logsin <= 24'd01419642;
                12'd2926: logsin <= 24'd01420511;
                12'd2927: logsin <= 24'd01421381;
                12'd2928: logsin <= 24'd01422250;
                12'd2929: logsin <= 24'd01423120;
                12'd2930: logsin <= 24'd01423989;
                12'd2931: logsin <= 24'd01424859;
                12'd2932: logsin <= 24'd01425728;
                12'd2933: logsin <= 24'd01426597;
                12'd2934: logsin <= 24'd01427467;
                12'd2935: logsin <= 24'd01428336;
                12'd2936: logsin <= 24'd01429205;
                12'd2937: logsin <= 24'd01430074;
                12'd2938: logsin <= 24'd01430943;
                12'd2939: logsin <= 24'd01431813;
                12'd2940: logsin <= 24'd01432682;
                12'd2941: logsin <= 24'd01433551;
                12'd2942: logsin <= 24'd01434420;
                12'd2943: logsin <= 24'd01435288;
                12'd2944: logsin <= 24'd01436157;
                12'd2945: logsin <= 24'd01437026;
                12'd2946: logsin <= 24'd01437895;
                12'd2947: logsin <= 24'd01438764;
                12'd2948: logsin <= 24'd01439632;
                12'd2949: logsin <= 24'd01440501;
                12'd2950: logsin <= 24'd01441370;
                12'd2951: logsin <= 24'd01442238;
                12'd2952: logsin <= 24'd01443106;
                12'd2953: logsin <= 24'd01443975;
                12'd2954: logsin <= 24'd01444843;
                12'd2955: logsin <= 24'd01445712;
                12'd2956: logsin <= 24'd01446580;
                12'd2957: logsin <= 24'd01447448;
                12'd2958: logsin <= 24'd01448316;
                12'd2959: logsin <= 24'd01449184;
                12'd2960: logsin <= 24'd01450052;
                12'd2961: logsin <= 24'd01450920;
                12'd2962: logsin <= 24'd01451788;
                12'd2963: logsin <= 24'd01452656;
                12'd2964: logsin <= 24'd01453523;
                12'd2965: logsin <= 24'd01454391;
                12'd2966: logsin <= 24'd01455259;
                12'd2967: logsin <= 24'd01456126;
                12'd2968: logsin <= 24'd01456994;
                12'd2969: logsin <= 24'd01457861;
                12'd2970: logsin <= 24'd01458728;
                12'd2971: logsin <= 24'd01459596;
                12'd2972: logsin <= 24'd01460463;
                12'd2973: logsin <= 24'd01461330;
                12'd2974: logsin <= 24'd01462197;
                12'd2975: logsin <= 24'd01463064;
                12'd2976: logsin <= 24'd01463931;
                12'd2977: logsin <= 24'd01464798;
                12'd2978: logsin <= 24'd01465664;
                12'd2979: logsin <= 24'd01466531;
                12'd2980: logsin <= 24'd01467398;
                12'd2981: logsin <= 24'd01468264;
                12'd2982: logsin <= 24'd01469130;
                12'd2983: logsin <= 24'd01469997;
                12'd2984: logsin <= 24'd01470863;
                12'd2985: logsin <= 24'd01471729;
                12'd2986: logsin <= 24'd01472595;
                12'd2987: logsin <= 24'd01473461;
                12'd2988: logsin <= 24'd01474327;
                12'd2989: logsin <= 24'd01475193;
                12'd2990: logsin <= 24'd01476059;
                12'd2991: logsin <= 24'd01476924;
                12'd2992: logsin <= 24'd01477790;
                12'd2993: logsin <= 24'd01478655;
                12'd2994: logsin <= 24'd01479521;
                12'd2995: logsin <= 24'd01480386;
                12'd2996: logsin <= 24'd01481251;
                12'd2997: logsin <= 24'd01482116;
                12'd2998: logsin <= 24'd01482981;
                12'd2999: logsin <= 24'd01483846;
                12'd3000: logsin <= 24'd01484711;
                12'd3001: logsin <= 24'd01485575;
                12'd3002: logsin <= 24'd01486440;
                12'd3003: logsin <= 24'd01487304;
                12'd3004: logsin <= 24'd01488169;
                12'd3005: logsin <= 24'd01489033;
                12'd3006: logsin <= 24'd01489897;
                12'd3007: logsin <= 24'd01490761;
                12'd3008: logsin <= 24'd01491625;
                12'd3009: logsin <= 24'd01492489;
                12'd3010: logsin <= 24'd01493353;
                12'd3011: logsin <= 24'd01494216;
                12'd3012: logsin <= 24'd01495080;
                12'd3013: logsin <= 24'd01495943;
                12'd3014: logsin <= 24'd01496806;
                12'd3015: logsin <= 24'd01497670;
                12'd3016: logsin <= 24'd01498533;
                12'd3017: logsin <= 24'd01499396;
                12'd3018: logsin <= 24'd01500258;
                12'd3019: logsin <= 24'd01501121;
                12'd3020: logsin <= 24'd01501984;
                12'd3021: logsin <= 24'd01502846;
                12'd3022: logsin <= 24'd01503708;
                12'd3023: logsin <= 24'd01504571;
                12'd3024: logsin <= 24'd01505433;
                12'd3025: logsin <= 24'd01506295;
                12'd3026: logsin <= 24'd01507157;
                12'd3027: logsin <= 24'd01508018;
                12'd3028: logsin <= 24'd01508880;
                12'd3029: logsin <= 24'd01509741;
                12'd3030: logsin <= 24'd01510603;
                12'd3031: logsin <= 24'd01511464;
                12'd3032: logsin <= 24'd01512325;
                12'd3033: logsin <= 24'd01513186;
                12'd3034: logsin <= 24'd01514047;
                12'd3035: logsin <= 24'd01514908;
                12'd3036: logsin <= 24'd01515768;
                12'd3037: logsin <= 24'd01516628;
                12'd3038: logsin <= 24'd01517489;
                12'd3039: logsin <= 24'd01518349;
                12'd3040: logsin <= 24'd01519209;
                12'd3041: logsin <= 24'd01520069;
                12'd3042: logsin <= 24'd01520929;
                12'd3043: logsin <= 24'd01521788;
                12'd3044: logsin <= 24'd01522648;
                12'd3045: logsin <= 24'd01523507;
                12'd3046: logsin <= 24'd01524366;
                12'd3047: logsin <= 24'd01525225;
                12'd3048: logsin <= 24'd01526084;
                12'd3049: logsin <= 24'd01526943;
                12'd3050: logsin <= 24'd01527801;
                12'd3051: logsin <= 24'd01528660;
                12'd3052: logsin <= 24'd01529518;
                12'd3053: logsin <= 24'd01530376;
                12'd3054: logsin <= 24'd01531234;
                12'd3055: logsin <= 24'd01532092;
                12'd3056: logsin <= 24'd01532949;
                12'd3057: logsin <= 24'd01533807;
                12'd3058: logsin <= 24'd01534664;
                12'd3059: logsin <= 24'd01535521;
                12'd3060: logsin <= 24'd01536378;
                12'd3061: logsin <= 24'd01537235;
                12'd3062: logsin <= 24'd01538092;
                12'd3063: logsin <= 24'd01538948;
                12'd3064: logsin <= 24'd01539805;
                12'd3065: logsin <= 24'd01540661;
                12'd3066: logsin <= 24'd01541517;
                12'd3067: logsin <= 24'd01542373;
                12'd3068: logsin <= 24'd01543229;
                12'd3069: logsin <= 24'd01544084;
                12'd3070: logsin <= 24'd01544939;
                12'd3071: logsin <= 24'd01545795;
                12'd3072: logsin <= 24'd01546650;
                12'd3073: logsin <= 24'd01547505;
                12'd3074: logsin <= 24'd01548359;
                12'd3075: logsin <= 24'd01549214;
                12'd3076: logsin <= 24'd01550068;
                12'd3077: logsin <= 24'd01550922;
                12'd3078: logsin <= 24'd01551776;
                12'd3079: logsin <= 24'd01552630;
                12'd3080: logsin <= 24'd01553484;
                12'd3081: logsin <= 24'd01554337;
                12'd3082: logsin <= 24'd01555190;
                12'd3083: logsin <= 24'd01556043;
                12'd3084: logsin <= 24'd01556896;
                12'd3085: logsin <= 24'd01557749;
                12'd3086: logsin <= 24'd01558601;
                12'd3087: logsin <= 24'd01559454;
                12'd3088: logsin <= 24'd01560306;
                12'd3089: logsin <= 24'd01561158;
                12'd3090: logsin <= 24'd01562009;
                12'd3091: logsin <= 24'd01562861;
                12'd3092: logsin <= 24'd01563712;
                12'd3093: logsin <= 24'd01564564;
                12'd3094: logsin <= 24'd01565414;
                12'd3095: logsin <= 24'd01566265;
                12'd3096: logsin <= 24'd01567116;
                12'd3097: logsin <= 24'd01567966;
                12'd3098: logsin <= 24'd01568816;
                12'd3099: logsin <= 24'd01569666;
                12'd3100: logsin <= 24'd01570516;
                12'd3101: logsin <= 24'd01571366;
                12'd3102: logsin <= 24'd01572215;
                12'd3103: logsin <= 24'd01573064;
                12'd3104: logsin <= 24'd01573913;
                12'd3105: logsin <= 24'd01574762;
                12'd3106: logsin <= 24'd01575610;
                12'd3107: logsin <= 24'd01576459;
                12'd3108: logsin <= 24'd01577307;
                12'd3109: logsin <= 24'd01578155;
                12'd3110: logsin <= 24'd01579002;
                12'd3111: logsin <= 24'd01579850;
                12'd3112: logsin <= 24'd01580697;
                12'd3113: logsin <= 24'd01581544;
                12'd3114: logsin <= 24'd01582391;
                12'd3115: logsin <= 24'd01583238;
                12'd3116: logsin <= 24'd01584084;
                12'd3117: logsin <= 24'd01584930;
                12'd3118: logsin <= 24'd01585776;
                12'd3119: logsin <= 24'd01586622;
                12'd3120: logsin <= 24'd01587467;
                12'd3121: logsin <= 24'd01588312;
                12'd3122: logsin <= 24'd01589157;
                12'd3123: logsin <= 24'd01590002;
                12'd3124: logsin <= 24'd01590847;
                12'd3125: logsin <= 24'd01591691;
                12'd3126: logsin <= 24'd01592535;
                12'd3127: logsin <= 24'd01593379;
                12'd3128: logsin <= 24'd01594223;
                12'd3129: logsin <= 24'd01595066;
                12'd3130: logsin <= 24'd01595909;
                12'd3131: logsin <= 24'd01596752;
                12'd3132: logsin <= 24'd01597595;
                12'd3133: logsin <= 24'd01598437;
                12'd3134: logsin <= 24'd01599280;
                12'd3135: logsin <= 24'd01600122;
                12'd3136: logsin <= 24'd01600963;
                12'd3137: logsin <= 24'd01601805;
                12'd3138: logsin <= 24'd01602646;
                12'd3139: logsin <= 24'd01603487;
                12'd3140: logsin <= 24'd01604328;
                12'd3141: logsin <= 24'd01605168;
                12'd3142: logsin <= 24'd01606009;
                12'd3143: logsin <= 24'd01606849;
                12'd3144: logsin <= 24'd01607688;
                12'd3145: logsin <= 24'd01608528;
                12'd3146: logsin <= 24'd01609367;
                12'd3147: logsin <= 24'd01610206;
                12'd3148: logsin <= 24'd01611045;
                12'd3149: logsin <= 24'd01611883;
                12'd3150: logsin <= 24'd01612721;
                12'd3151: logsin <= 24'd01613559;
                12'd3152: logsin <= 24'd01614397;
                12'd3153: logsin <= 24'd01615234;
                12'd3154: logsin <= 24'd01616071;
                12'd3155: logsin <= 24'd01616908;
                12'd3156: logsin <= 24'd01617745;
                12'd3157: logsin <= 24'd01618581;
                12'd3158: logsin <= 24'd01619417;
                12'd3159: logsin <= 24'd01620253;
                12'd3160: logsin <= 24'd01621089;
                12'd3161: logsin <= 24'd01621924;
                12'd3162: logsin <= 24'd01622759;
                12'd3163: logsin <= 24'd01623594;
                12'd3164: logsin <= 24'd01624428;
                12'd3165: logsin <= 24'd01625262;
                12'd3166: logsin <= 24'd01626096;
                12'd3167: logsin <= 24'd01626930;
                12'd3168: logsin <= 24'd01627763;
                12'd3169: logsin <= 24'd01628596;
                12'd3170: logsin <= 24'd01629429;
                12'd3171: logsin <= 24'd01630261;
                12'd3172: logsin <= 24'd01631094;
                12'd3173: logsin <= 24'd01631925;
                12'd3174: logsin <= 24'd01632757;
                12'd3175: logsin <= 24'd01633588;
                12'd3176: logsin <= 24'd01634419;
                12'd3177: logsin <= 24'd01635250;
                12'd3178: logsin <= 24'd01636081;
                12'd3179: logsin <= 24'd01636911;
                12'd3180: logsin <= 24'd01637740;
                12'd3181: logsin <= 24'd01638570;
                12'd3182: logsin <= 24'd01639399;
                12'd3183: logsin <= 24'd01640228;
                12'd3184: logsin <= 24'd01641057;
                12'd3185: logsin <= 24'd01641885;
                12'd3186: logsin <= 24'd01642713;
                12'd3187: logsin <= 24'd01643541;
                12'd3188: logsin <= 24'd01644368;
                12'd3189: logsin <= 24'd01645196;
                12'd3190: logsin <= 24'd01646022;
                12'd3191: logsin <= 24'd01646849;
                12'd3192: logsin <= 24'd01647675;
                12'd3193: logsin <= 24'd01648501;
                12'd3194: logsin <= 24'd01649327;
                12'd3195: logsin <= 24'd01650152;
                12'd3196: logsin <= 24'd01650977;
                12'd3197: logsin <= 24'd01651801;
                12'd3198: logsin <= 24'd01652626;
                12'd3199: logsin <= 24'd01653450;
                12'd3200: logsin <= 24'd01654273;
                12'd3201: logsin <= 24'd01655097;
                12'd3202: logsin <= 24'd01655920;
                12'd3203: logsin <= 24'd01656742;
                12'd3204: logsin <= 24'd01657565;
                12'd3205: logsin <= 24'd01658387;
                12'd3206: logsin <= 24'd01659209;
                12'd3207: logsin <= 24'd01660030;
                12'd3208: logsin <= 24'd01660851;
                12'd3209: logsin <= 24'd01661672;
                12'd3210: logsin <= 24'd01662492;
                12'd3211: logsin <= 24'd01663312;
                12'd3212: logsin <= 24'd01664132;
                12'd3213: logsin <= 24'd01664951;
                12'd3214: logsin <= 24'd01665770;
                12'd3215: logsin <= 24'd01666589;
                12'd3216: logsin <= 24'd01667407;
                12'd3217: logsin <= 24'd01668225;
                12'd3218: logsin <= 24'd01669043;
                12'd3219: logsin <= 24'd01669860;
                12'd3220: logsin <= 24'd01670677;
                12'd3221: logsin <= 24'd01671494;
                12'd3222: logsin <= 24'd01672310;
                12'd3223: logsin <= 24'd01673126;
                12'd3224: logsin <= 24'd01673942;
                12'd3225: logsin <= 24'd01674757;
                12'd3226: logsin <= 24'd01675572;
                12'd3227: logsin <= 24'd01676387;
                12'd3228: logsin <= 24'd01677201;
                12'd3229: logsin <= 24'd01678015;
                12'd3230: logsin <= 24'd01678828;
                12'd3231: logsin <= 24'd01679641;
                12'd3232: logsin <= 24'd01680454;
                12'd3233: logsin <= 24'd01681266;
                12'd3234: logsin <= 24'd01682078;
                12'd3235: logsin <= 24'd01682890;
                12'd3236: logsin <= 24'd01683701;
                12'd3237: logsin <= 24'd01684512;
                12'd3238: logsin <= 24'd01685323;
                12'd3239: logsin <= 24'd01686133;
                12'd3240: logsin <= 24'd01686943;
                12'd3241: logsin <= 24'd01687752;
                12'd3242: logsin <= 24'd01688561;
                12'd3243: logsin <= 24'd01689370;
                12'd3244: logsin <= 24'd01690178;
                12'd3245: logsin <= 24'd01690986;
                12'd3246: logsin <= 24'd01691794;
                12'd3247: logsin <= 24'd01692601;
                12'd3248: logsin <= 24'd01693407;
                12'd3249: logsin <= 24'd01694214;
                12'd3250: logsin <= 24'd01695020;
                12'd3251: logsin <= 24'd01695825;
                12'd3252: logsin <= 24'd01696631;
                12'd3253: logsin <= 24'd01697436;
                12'd3254: logsin <= 24'd01698240;
                12'd3255: logsin <= 24'd01699044;
                12'd3256: logsin <= 24'd01699848;
                12'd3257: logsin <= 24'd01700651;
                12'd3258: logsin <= 24'd01701454;
                12'd3259: logsin <= 24'd01702256;
                12'd3260: logsin <= 24'd01703058;
                12'd3261: logsin <= 24'd01703860;
                12'd3262: logsin <= 24'd01704661;
                12'd3263: logsin <= 24'd01705462;
                12'd3264: logsin <= 24'd01706263;
                12'd3265: logsin <= 24'd01707063;
                12'd3266: logsin <= 24'd01707863;
                12'd3267: logsin <= 24'd01708662;
                12'd3268: logsin <= 24'd01709461;
                12'd3269: logsin <= 24'd01710259;
                12'd3270: logsin <= 24'd01711057;
                12'd3271: logsin <= 24'd01711855;
                12'd3272: logsin <= 24'd01712652;
                12'd3273: logsin <= 24'd01713449;
                12'd3274: logsin <= 24'd01714245;
                12'd3275: logsin <= 24'd01715041;
                12'd3276: logsin <= 24'd01715837;
                12'd3277: logsin <= 24'd01716632;
                12'd3278: logsin <= 24'd01717426;
                12'd3279: logsin <= 24'd01718221;
                12'd3280: logsin <= 24'd01719014;
                12'd3281: logsin <= 24'd01719808;
                12'd3282: logsin <= 24'd01720601;
                12'd3283: logsin <= 24'd01721393;
                12'd3284: logsin <= 24'd01722186;
                12'd3285: logsin <= 24'd01722977;
                12'd3286: logsin <= 24'd01723768;
                12'd3287: logsin <= 24'd01724559;
                12'd3288: logsin <= 24'd01725350;
                12'd3289: logsin <= 24'd01726140;
                12'd3290: logsin <= 24'd01726929;
                12'd3291: logsin <= 24'd01727718;
                12'd3292: logsin <= 24'd01728507;
                12'd3293: logsin <= 24'd01729295;
                12'd3294: logsin <= 24'd01730083;
                12'd3295: logsin <= 24'd01730870;
                12'd3296: logsin <= 24'd01731657;
                12'd3297: logsin <= 24'd01732443;
                12'd3298: logsin <= 24'd01733229;
                12'd3299: logsin <= 24'd01734015;
                12'd3300: logsin <= 24'd01734800;
                12'd3301: logsin <= 24'd01735584;
                12'd3302: logsin <= 24'd01736369;
                12'd3303: logsin <= 24'd01737152;
                12'd3304: logsin <= 24'd01737936;
                12'd3305: logsin <= 24'd01738718;
                12'd3306: logsin <= 24'd01739501;
                12'd3307: logsin <= 24'd01740282;
                12'd3308: logsin <= 24'd01741064;
                12'd3309: logsin <= 24'd01741845;
                12'd3310: logsin <= 24'd01742625;
                12'd3311: logsin <= 24'd01743405;
                12'd3312: logsin <= 24'd01744185;
                12'd3313: logsin <= 24'd01744964;
                12'd3314: logsin <= 24'd01745742;
                12'd3315: logsin <= 24'd01746520;
                12'd3316: logsin <= 24'd01747298;
                12'd3317: logsin <= 24'd01748075;
                12'd3318: logsin <= 24'd01748852;
                12'd3319: logsin <= 24'd01749628;
                12'd3320: logsin <= 24'd01750404;
                12'd3321: logsin <= 24'd01751179;
                12'd3322: logsin <= 24'd01751954;
                12'd3323: logsin <= 24'd01752728;
                12'd3324: logsin <= 24'd01753502;
                12'd3325: logsin <= 24'd01754275;
                12'd3326: logsin <= 24'd01755048;
                12'd3327: logsin <= 24'd01755820;
                12'd3328: logsin <= 24'd01756592;
                12'd3329: logsin <= 24'd01757363;
                12'd3330: logsin <= 24'd01758134;
                12'd3331: logsin <= 24'd01758904;
                12'd3332: logsin <= 24'd01759674;
                12'd3333: logsin <= 24'd01760444;
                12'd3334: logsin <= 24'd01761212;
                12'd3335: logsin <= 24'd01761981;
                12'd3336: logsin <= 24'd01762749;
                12'd3337: logsin <= 24'd01763516;
                12'd3338: logsin <= 24'd01764283;
                12'd3339: logsin <= 24'd01765049;
                12'd3340: logsin <= 24'd01765815;
                12'd3341: logsin <= 24'd01766580;
                12'd3342: logsin <= 24'd01767345;
                12'd3343: logsin <= 24'd01768109;
                12'd3344: logsin <= 24'd01768873;
                12'd3345: logsin <= 24'd01769636;
                12'd3346: logsin <= 24'd01770399;
                12'd3347: logsin <= 24'd01771161;
                12'd3348: logsin <= 24'd01771923;
                12'd3349: logsin <= 24'd01772684;
                12'd3350: logsin <= 24'd01773445;
                12'd3351: logsin <= 24'd01774205;
                12'd3352: logsin <= 24'd01774964;
                12'd3353: logsin <= 24'd01775723;
                12'd3354: logsin <= 24'd01776482;
                12'd3355: logsin <= 24'd01777240;
                12'd3356: logsin <= 24'd01777998;
                12'd3357: logsin <= 24'd01778754;
                12'd3358: logsin <= 24'd01779511;
                12'd3359: logsin <= 24'd01780267;
                12'd3360: logsin <= 24'd01781022;
                12'd3361: logsin <= 24'd01781777;
                12'd3362: logsin <= 24'd01782531;
                12'd3363: logsin <= 24'd01783285;
                12'd3364: logsin <= 24'd01784038;
                12'd3365: logsin <= 24'd01784791;
                12'd3366: logsin <= 24'd01785543;
                12'd3367: logsin <= 24'd01786294;
                12'd3368: logsin <= 24'd01787045;
                12'd3369: logsin <= 24'd01787796;
                12'd3370: logsin <= 24'd01788546;
                12'd3371: logsin <= 24'd01789295;
                12'd3372: logsin <= 24'd01790044;
                12'd3373: logsin <= 24'd01790792;
                12'd3374: logsin <= 24'd01791540;
                12'd3375: logsin <= 24'd01792287;
                12'd3376: logsin <= 24'd01793033;
                12'd3377: logsin <= 24'd01793779;
                12'd3378: logsin <= 24'd01794525;
                12'd3379: logsin <= 24'd01795270;
                12'd3380: logsin <= 24'd01796014;
                12'd3381: logsin <= 24'd01796758;
                12'd3382: logsin <= 24'd01797501;
                12'd3383: logsin <= 24'd01798243;
                12'd3384: logsin <= 24'd01798985;
                12'd3385: logsin <= 24'd01799727;
                12'd3386: logsin <= 24'd01800468;
                12'd3387: logsin <= 24'd01801208;
                12'd3388: logsin <= 24'd01801948;
                12'd3389: logsin <= 24'd01802687;
                12'd3390: logsin <= 24'd01803425;
                12'd3391: logsin <= 24'd01804163;
                12'd3392: logsin <= 24'd01804901;
                12'd3393: logsin <= 24'd01805638;
                12'd3394: logsin <= 24'd01806374;
                12'd3395: logsin <= 24'd01807109;
                12'd3396: logsin <= 24'd01807845;
                12'd3397: logsin <= 24'd01808579;
                12'd3398: logsin <= 24'd01809313;
                12'd3399: logsin <= 24'd01810046;
                12'd3400: logsin <= 24'd01810779;
                12'd3401: logsin <= 24'd01811511;
                12'd3402: logsin <= 24'd01812242;
                12'd3403: logsin <= 24'd01812973;
                12'd3404: logsin <= 24'd01813704;
                12'd3405: logsin <= 24'd01814433;
                12'd3406: logsin <= 24'd01815162;
                12'd3407: logsin <= 24'd01815891;
                12'd3408: logsin <= 24'd01816619;
                12'd3409: logsin <= 24'd01817346;
                12'd3410: logsin <= 24'd01818072;
                12'd3411: logsin <= 24'd01818798;
                12'd3412: logsin <= 24'd01819524;
                12'd3413: logsin <= 24'd01820249;
                12'd3414: logsin <= 24'd01820973;
                12'd3415: logsin <= 24'd01821696;
                12'd3416: logsin <= 24'd01822419;
                12'd3417: logsin <= 24'd01823142;
                12'd3418: logsin <= 24'd01823863;
                12'd3419: logsin <= 24'd01824585;
                12'd3420: logsin <= 24'd01825305;
                12'd3421: logsin <= 24'd01826025;
                12'd3422: logsin <= 24'd01826744;
                12'd3423: logsin <= 24'd01827463;
                12'd3424: logsin <= 24'd01828181;
                12'd3425: logsin <= 24'd01828898;
                12'd3426: logsin <= 24'd01829615;
                12'd3427: logsin <= 24'd01830331;
                12'd3428: logsin <= 24'd01831046;
                12'd3429: logsin <= 24'd01831761;
                12'd3430: logsin <= 24'd01832475;
                12'd3431: logsin <= 24'd01833188;
                12'd3432: logsin <= 24'd01833901;
                12'd3433: logsin <= 24'd01834613;
                12'd3434: logsin <= 24'd01835325;
                12'd3435: logsin <= 24'd01836036;
                12'd3436: logsin <= 24'd01836746;
                12'd3437: logsin <= 24'd01837456;
                12'd3438: logsin <= 24'd01838165;
                12'd3439: logsin <= 24'd01838873;
                12'd3440: logsin <= 24'd01839581;
                12'd3441: logsin <= 24'd01840288;
                12'd3442: logsin <= 24'd01840994;
                12'd3443: logsin <= 24'd01841700;
                12'd3444: logsin <= 24'd01842405;
                12'd3445: logsin <= 24'd01843109;
                12'd3446: logsin <= 24'd01843813;
                12'd3447: logsin <= 24'd01844516;
                12'd3448: logsin <= 24'd01845218;
                12'd3449: logsin <= 24'd01845920;
                12'd3450: logsin <= 24'd01846621;
                12'd3451: logsin <= 24'd01847321;
                12'd3452: logsin <= 24'd01848021;
                12'd3453: logsin <= 24'd01848720;
                12'd3454: logsin <= 24'd01849418;
                12'd3455: logsin <= 24'd01850116;
                12'd3456: logsin <= 24'd01850813;
                12'd3457: logsin <= 24'd01851509;
                12'd3458: logsin <= 24'd01852205;
                12'd3459: logsin <= 24'd01852900;
                12'd3460: logsin <= 24'd01853594;
                12'd3461: logsin <= 24'd01854288;
                12'd3462: logsin <= 24'd01854981;
                12'd3463: logsin <= 24'd01855673;
                12'd3464: logsin <= 24'd01856364;
                12'd3465: logsin <= 24'd01857055;
                12'd3466: logsin <= 24'd01857745;
                12'd3467: logsin <= 24'd01858435;
                12'd3468: logsin <= 24'd01859123;
                12'd3469: logsin <= 24'd01859811;
                12'd3470: logsin <= 24'd01860499;
                12'd3471: logsin <= 24'd01861185;
                12'd3472: logsin <= 24'd01861871;
                12'd3473: logsin <= 24'd01862557;
                12'd3474: logsin <= 24'd01863241;
                12'd3475: logsin <= 24'd01863925;
                12'd3476: logsin <= 24'd01864608;
                12'd3477: logsin <= 24'd01865290;
                12'd3478: logsin <= 24'd01865972;
                12'd3479: logsin <= 24'd01866653;
                12'd3480: logsin <= 24'd01867333;
                12'd3481: logsin <= 24'd01868013;
                12'd3482: logsin <= 24'd01868692;
                12'd3483: logsin <= 24'd01869370;
                12'd3484: logsin <= 24'd01870047;
                12'd3485: logsin <= 24'd01870724;
                12'd3486: logsin <= 24'd01871400;
                12'd3487: logsin <= 24'd01872075;
                12'd3488: logsin <= 24'd01872749;
                12'd3489: logsin <= 24'd01873423;
                12'd3490: logsin <= 24'd01874096;
                12'd3491: logsin <= 24'd01874768;
                12'd3492: logsin <= 24'd01875440;
                12'd3493: logsin <= 24'd01876111;
                12'd3494: logsin <= 24'd01876781;
                12'd3495: logsin <= 24'd01877450;
                12'd3496: logsin <= 24'd01878119;
                12'd3497: logsin <= 24'd01878787;
                12'd3498: logsin <= 24'd01879454;
                12'd3499: logsin <= 24'd01880120;
                12'd3500: logsin <= 24'd01880786;
                12'd3501: logsin <= 24'd01881451;
                12'd3502: logsin <= 24'd01882115;
                12'd3503: logsin <= 24'd01882779;
                12'd3504: logsin <= 24'd01883441;
                12'd3505: logsin <= 24'd01884103;
                12'd3506: logsin <= 24'd01884764;
                12'd3507: logsin <= 24'd01885425;
                12'd3508: logsin <= 24'd01886084;
                12'd3509: logsin <= 24'd01886743;
                12'd3510: logsin <= 24'd01887401;
                12'd3511: logsin <= 24'd01888059;
                12'd3512: logsin <= 24'd01888715;
                12'd3513: logsin <= 24'd01889371;
                12'd3514: logsin <= 24'd01890026;
                12'd3515: logsin <= 24'd01890681;
                12'd3516: logsin <= 24'd01891334;
                12'd3517: logsin <= 24'd01891987;
                12'd3518: logsin <= 24'd01892639;
                12'd3519: logsin <= 24'd01893290;
                12'd3520: logsin <= 24'd01893941;
                12'd3521: logsin <= 24'd01894590;
                12'd3522: logsin <= 24'd01895239;
                12'd3523: logsin <= 24'd01895887;
                12'd3524: logsin <= 24'd01896535;
                12'd3525: logsin <= 24'd01897181;
                12'd3526: logsin <= 24'd01897827;
                12'd3527: logsin <= 24'd01898472;
                12'd3528: logsin <= 24'd01899116;
                12'd3529: logsin <= 24'd01899759;
                12'd3530: logsin <= 24'd01900402;
                12'd3531: logsin <= 24'd01901044;
                12'd3532: logsin <= 24'd01901685;
                12'd3533: logsin <= 24'd01902325;
                12'd3534: logsin <= 24'd01902965;
                12'd3535: logsin <= 24'd01903603;
                12'd3536: logsin <= 24'd01904241;
                12'd3537: logsin <= 24'd01904878;
                12'd3538: logsin <= 24'd01905515;
                12'd3539: logsin <= 24'd01906150;
                12'd3540: logsin <= 24'd01906785;
                12'd3541: logsin <= 24'd01907418;
                12'd3542: logsin <= 24'd01908052;
                12'd3543: logsin <= 24'd01908684;
                12'd3544: logsin <= 24'd01909315;
                12'd3545: logsin <= 24'd01909946;
                12'd3546: logsin <= 24'd01910576;
                12'd3547: logsin <= 24'd01911205;
                12'd3548: logsin <= 24'd01911833;
                12'd3549: logsin <= 24'd01912460;
                12'd3550: logsin <= 24'd01913087;
                12'd3551: logsin <= 24'd01913712;
                12'd3552: logsin <= 24'd01914337;
                12'd3553: logsin <= 24'd01914961;
                12'd3554: logsin <= 24'd01915584;
                12'd3555: logsin <= 24'd01916207;
                12'd3556: logsin <= 24'd01916828;
                12'd3557: logsin <= 24'd01917449;
                12'd3558: logsin <= 24'd01918069;
                12'd3559: logsin <= 24'd01918688;
                12'd3560: logsin <= 24'd01919306;
                12'd3561: logsin <= 24'd01919924;
                12'd3562: logsin <= 24'd01920540;
                12'd3563: logsin <= 24'd01921156;
                12'd3564: logsin <= 24'd01921771;
                12'd3565: logsin <= 24'd01922385;
                12'd3566: logsin <= 24'd01922998;
                12'd3567: logsin <= 24'd01923611;
                12'd3568: logsin <= 24'd01924222;
                12'd3569: logsin <= 24'd01924833;
                12'd3570: logsin <= 24'd01925443;
                12'd3571: logsin <= 24'd01926052;
                12'd3572: logsin <= 24'd01926660;
                12'd3573: logsin <= 24'd01927267;
                12'd3574: logsin <= 24'd01927873;
                12'd3575: logsin <= 24'd01928479;
                12'd3576: logsin <= 24'd01929084;
                12'd3577: logsin <= 24'd01929687;
                12'd3578: logsin <= 24'd01930290;
                12'd3579: logsin <= 24'd01930893;
                12'd3580: logsin <= 24'd01931494;
                12'd3581: logsin <= 24'd01932094;
                12'd3582: logsin <= 24'd01932694;
                12'd3583: logsin <= 24'd01933292;
                12'd3584: logsin <= 24'd01933890;
                12'd3585: logsin <= 24'd01934487;
                12'd3586: logsin <= 24'd01935083;
                12'd3587: logsin <= 24'd01935678;
                12'd3588: logsin <= 24'd01936273;
                12'd3589: logsin <= 24'd01936866;
                12'd3590: logsin <= 24'd01937458;
                12'd3591: logsin <= 24'd01938050;
                12'd3592: logsin <= 24'd01938641;
                12'd3593: logsin <= 24'd01939231;
                12'd3594: logsin <= 24'd01939820;
                12'd3595: logsin <= 24'd01940408;
                12'd3596: logsin <= 24'd01940995;
                12'd3597: logsin <= 24'd01941581;
                12'd3598: logsin <= 24'd01942167;
                12'd3599: logsin <= 24'd01942751;
                12'd3600: logsin <= 24'd01943335;
                12'd3601: logsin <= 24'd01943918;
                12'd3602: logsin <= 24'd01944500;
                12'd3603: logsin <= 24'd01945081;
                12'd3604: logsin <= 24'd01945661;
                12'd3605: logsin <= 24'd01946240;
                12'd3606: logsin <= 24'd01946818;
                12'd3607: logsin <= 24'd01947396;
                12'd3608: logsin <= 24'd01947972;
                12'd3609: logsin <= 24'd01948548;
                12'd3610: logsin <= 24'd01949122;
                12'd3611: logsin <= 24'd01949696;
                12'd3612: logsin <= 24'd01950269;
                12'd3613: logsin <= 24'd01950841;
                12'd3614: logsin <= 24'd01951412;
                12'd3615: logsin <= 24'd01951982;
                12'd3616: logsin <= 24'd01952551;
                12'd3617: logsin <= 24'd01953119;
                12'd3618: logsin <= 24'd01953686;
                12'd3619: logsin <= 24'd01954253;
                12'd3620: logsin <= 24'd01954818;
                12'd3621: logsin <= 24'd01955383;
                12'd3622: logsin <= 24'd01955947;
                12'd3623: logsin <= 24'd01956509;
                12'd3624: logsin <= 24'd01957071;
                12'd3625: logsin <= 24'd01957632;
                12'd3626: logsin <= 24'd01958192;
                12'd3627: logsin <= 24'd01958751;
                12'd3628: logsin <= 24'd01959309;
                12'd3629: logsin <= 24'd01959866;
                12'd3630: logsin <= 24'd01960422;
                12'd3631: logsin <= 24'd01960977;
                12'd3632: logsin <= 24'd01961532;
                12'd3633: logsin <= 24'd01962085;
                12'd3634: logsin <= 24'd01962637;
                12'd3635: logsin <= 24'd01963189;
                12'd3636: logsin <= 24'd01963739;
                12'd3637: logsin <= 24'd01964289;
                12'd3638: logsin <= 24'd01964838;
                12'd3639: logsin <= 24'd01965385;
                12'd3640: logsin <= 24'd01965932;
                12'd3641: logsin <= 24'd01966478;
                12'd3642: logsin <= 24'd01967023;
                12'd3643: logsin <= 24'd01967566;
                12'd3644: logsin <= 24'd01968109;
                12'd3645: logsin <= 24'd01968651;
                12'd3646: logsin <= 24'd01969192;
                12'd3647: logsin <= 24'd01969732;
                12'd3648: logsin <= 24'd01970271;
                12'd3649: logsin <= 24'd01970810;
                12'd3650: logsin <= 24'd01971347;
                12'd3651: logsin <= 24'd01971883;
                12'd3652: logsin <= 24'd01972418;
                12'd3653: logsin <= 24'd01972952;
                12'd3654: logsin <= 24'd01973485;
                12'd3655: logsin <= 24'd01974018;
                12'd3656: logsin <= 24'd01974549;
                12'd3657: logsin <= 24'd01975079;
                12'd3658: logsin <= 24'd01975609;
                12'd3659: logsin <= 24'd01976137;
                12'd3660: logsin <= 24'd01976665;
                12'd3661: logsin <= 24'd01977191;
                12'd3662: logsin <= 24'd01977716;
                12'd3663: logsin <= 24'd01978241;
                12'd3664: logsin <= 24'd01978764;
                12'd3665: logsin <= 24'd01979287;
                12'd3666: logsin <= 24'd01979808;
                12'd3667: logsin <= 24'd01980329;
                12'd3668: logsin <= 24'd01980848;
                12'd3669: logsin <= 24'd01981367;
                12'd3670: logsin <= 24'd01981884;
                12'd3671: logsin <= 24'd01982401;
                12'd3672: logsin <= 24'd01982916;
                12'd3673: logsin <= 24'd01983431;
                12'd3674: logsin <= 24'd01983945;
                12'd3675: logsin <= 24'd01984457;
                12'd3676: logsin <= 24'd01984969;
                12'd3677: logsin <= 24'd01985479;
                12'd3678: logsin <= 24'd01985989;
                12'd3679: logsin <= 24'd01986497;
                12'd3680: logsin <= 24'd01987005;
                12'd3681: logsin <= 24'd01987511;
                12'd3682: logsin <= 24'd01988017;
                12'd3683: logsin <= 24'd01988521;
                12'd3684: logsin <= 24'd01989025;
                12'd3685: logsin <= 24'd01989527;
                12'd3686: logsin <= 24'd01990029;
                12'd3687: logsin <= 24'd01990529;
                12'd3688: logsin <= 24'd01991028;
                12'd3689: logsin <= 24'd01991527;
                12'd3690: logsin <= 24'd01992024;
                12'd3691: logsin <= 24'd01992521;
                12'd3692: logsin <= 24'd01993016;
                12'd3693: logsin <= 24'd01993510;
                12'd3694: logsin <= 24'd01994003;
                12'd3695: logsin <= 24'd01994496;
                12'd3696: logsin <= 24'd01994987;
                12'd3697: logsin <= 24'd01995477;
                12'd3698: logsin <= 24'd01995966;
                12'd3699: logsin <= 24'd01996454;
                12'd3700: logsin <= 24'd01996941;
                12'd3701: logsin <= 24'd01997427;
                12'd3702: logsin <= 24'd01997912;
                12'd3703: logsin <= 24'd01998396;
                12'd3704: logsin <= 24'd01998879;
                12'd3705: logsin <= 24'd01999361;
                12'd3706: logsin <= 24'd01999842;
                12'd3707: logsin <= 24'd02000322;
                12'd3708: logsin <= 24'd02000801;
                12'd3709: logsin <= 24'd02001278;
                12'd3710: logsin <= 24'd02001755;
                12'd3711: logsin <= 24'd02002231;
                12'd3712: logsin <= 24'd02002705;
                12'd3713: logsin <= 24'd02003179;
                12'd3714: logsin <= 24'd02003651;
                12'd3715: logsin <= 24'd02004123;
                12'd3716: logsin <= 24'd02004593;
                12'd3717: logsin <= 24'd02005062;
                12'd3718: logsin <= 24'd02005531;
                12'd3719: logsin <= 24'd02005998;
                12'd3720: logsin <= 24'd02006464;
                12'd3721: logsin <= 24'd02006929;
                12'd3722: logsin <= 24'd02007393;
                12'd3723: logsin <= 24'd02007856;
                12'd3724: logsin <= 24'd02008318;
                12'd3725: logsin <= 24'd02008778;
                12'd3726: logsin <= 24'd02009238;
                12'd3727: logsin <= 24'd02009697;
                12'd3728: logsin <= 24'd02010154;
                12'd3729: logsin <= 24'd02010611;
                12'd3730: logsin <= 24'd02011066;
                12'd3731: logsin <= 24'd02011521;
                12'd3732: logsin <= 24'd02011974;
                12'd3733: logsin <= 24'd02012426;
                12'd3734: logsin <= 24'd02012877;
                12'd3735: logsin <= 24'd02013327;
                12'd3736: logsin <= 24'd02013776;
                12'd3737: logsin <= 24'd02014224;
                12'd3738: logsin <= 24'd02014671;
                12'd3739: logsin <= 24'd02015117;
                12'd3740: logsin <= 24'd02015561;
                12'd3741: logsin <= 24'd02016005;
                12'd3742: logsin <= 24'd02016447;
                12'd3743: logsin <= 24'd02016889;
                12'd3744: logsin <= 24'd02017329;
                12'd3745: logsin <= 24'd02017768;
                12'd3746: logsin <= 24'd02018206;
                12'd3747: logsin <= 24'd02018643;
                12'd3748: logsin <= 24'd02019079;
                12'd3749: logsin <= 24'd02019514;
                12'd3750: logsin <= 24'd02019948;
                12'd3751: logsin <= 24'd02020380;
                12'd3752: logsin <= 24'd02020812;
                12'd3753: logsin <= 24'd02021242;
                12'd3754: logsin <= 24'd02021671;
                12'd3755: logsin <= 24'd02022100;
                12'd3756: logsin <= 24'd02022527;
                12'd3757: logsin <= 24'd02022953;
                12'd3758: logsin <= 24'd02023378;
                12'd3759: logsin <= 24'd02023801;
                12'd3760: logsin <= 24'd02024224;
                12'd3761: logsin <= 24'd02024645;
                12'd3762: logsin <= 24'd02025066;
                12'd3763: logsin <= 24'd02025485;
                12'd3764: logsin <= 24'd02025903;
                12'd3765: logsin <= 24'd02026320;
                12'd3766: logsin <= 24'd02026736;
                12'd3767: logsin <= 24'd02027151;
                12'd3768: logsin <= 24'd02027565;
                12'd3769: logsin <= 24'd02027977;
                12'd3770: logsin <= 24'd02028389;
                12'd3771: logsin <= 24'd02028799;
                12'd3772: logsin <= 24'd02029208;
                12'd3773: logsin <= 24'd02029617;
                12'd3774: logsin <= 24'd02030024;
                12'd3775: logsin <= 24'd02030429;
                12'd3776: logsin <= 24'd02030834;
                12'd3777: logsin <= 24'd02031238;
                12'd3778: logsin <= 24'd02031640;
                12'd3779: logsin <= 24'd02032041;
                12'd3780: logsin <= 24'd02032442;
                12'd3781: logsin <= 24'd02032841;
                12'd3782: logsin <= 24'd02033238;
                12'd3783: logsin <= 24'd02033635;
                12'd3784: logsin <= 24'd02034031;
                12'd3785: logsin <= 24'd02034425;
                12'd3786: logsin <= 24'd02034819;
                12'd3787: logsin <= 24'd02035211;
                12'd3788: logsin <= 24'd02035602;
                12'd3789: logsin <= 24'd02035992;
                12'd3790: logsin <= 24'd02036380;
                12'd3791: logsin <= 24'd02036768;
                12'd3792: logsin <= 24'd02037155;
                12'd3793: logsin <= 24'd02037540;
                12'd3794: logsin <= 24'd02037924;
                12'd3795: logsin <= 24'd02038307;
                12'd3796: logsin <= 24'd02038689;
                12'd3797: logsin <= 24'd02039070;
                12'd3798: logsin <= 24'd02039449;
                12'd3799: logsin <= 24'd02039827;
                12'd3800: logsin <= 24'd02040205;
                12'd3801: logsin <= 24'd02040581;
                12'd3802: logsin <= 24'd02040956;
                12'd3803: logsin <= 24'd02041329;
                12'd3804: logsin <= 24'd02041702;
                12'd3805: logsin <= 24'd02042073;
                12'd3806: logsin <= 24'd02042444;
                12'd3807: logsin <= 24'd02042813;
                12'd3808: logsin <= 24'd02043181;
                12'd3809: logsin <= 24'd02043547;
                12'd3810: logsin <= 24'd02043913;
                12'd3811: logsin <= 24'd02044277;
                12'd3812: logsin <= 24'd02044641;
                12'd3813: logsin <= 24'd02045003;
                12'd3814: logsin <= 24'd02045364;
                12'd3815: logsin <= 24'd02045723;
                12'd3816: logsin <= 24'd02046082;
                12'd3817: logsin <= 24'd02046439;
                12'd3818: logsin <= 24'd02046795;
                12'd3819: logsin <= 24'd02047150;
                12'd3820: logsin <= 24'd02047504;
                12'd3821: logsin <= 24'd02047857;
                12'd3822: logsin <= 24'd02048208;
                12'd3823: logsin <= 24'd02048559;
                12'd3824: logsin <= 24'd02048908;
                12'd3825: logsin <= 24'd02049256;
                12'd3826: logsin <= 24'd02049602;
                12'd3827: logsin <= 24'd02049948;
                12'd3828: logsin <= 24'd02050292;
                12'd3829: logsin <= 24'd02050636;
                12'd3830: logsin <= 24'd02050978;
                12'd3831: logsin <= 24'd02051318;
                12'd3832: logsin <= 24'd02051658;
                12'd3833: logsin <= 24'd02051996;
                12'd3834: logsin <= 24'd02052334;
                12'd3835: logsin <= 24'd02052670;
                12'd3836: logsin <= 24'd02053004;
                12'd3837: logsin <= 24'd02053338;
                12'd3838: logsin <= 24'd02053670;
                12'd3839: logsin <= 24'd02054002;
                12'd3840: logsin <= 24'd02054332;
                12'd3841: logsin <= 24'd02054661;
                12'd3842: logsin <= 24'd02054988;
                12'd3843: logsin <= 24'd02055315;
                12'd3844: logsin <= 24'd02055640;
                12'd3845: logsin <= 24'd02055964;
                12'd3846: logsin <= 24'd02056287;
                12'd3847: logsin <= 24'd02056608;
                12'd3848: logsin <= 24'd02056929;
                12'd3849: logsin <= 24'd02057248;
                12'd3850: logsin <= 24'd02057566;
                12'd3851: logsin <= 24'd02057883;
                12'd3852: logsin <= 24'd02058198;
                12'd3853: logsin <= 24'd02058512;
                12'd3854: logsin <= 24'd02058826;
                12'd3855: logsin <= 24'd02059137;
                12'd3856: logsin <= 24'd02059448;
                12'd3857: logsin <= 24'd02059758;
                12'd3858: logsin <= 24'd02060066;
                12'd3859: logsin <= 24'd02060373;
                12'd3860: logsin <= 24'd02060679;
                12'd3861: logsin <= 24'd02060983;
                12'd3862: logsin <= 24'd02061287;
                12'd3863: logsin <= 24'd02061589;
                12'd3864: logsin <= 24'd02061890;
                12'd3865: logsin <= 24'd02062190;
                12'd3866: logsin <= 24'd02062488;
                12'd3867: logsin <= 24'd02062785;
                12'd3868: logsin <= 24'd02063081;
                12'd3869: logsin <= 24'd02063376;
                12'd3870: logsin <= 24'd02063670;
                12'd3871: logsin <= 24'd02063962;
                12'd3872: logsin <= 24'd02064253;
                12'd3873: logsin <= 24'd02064543;
                12'd3874: logsin <= 24'd02064832;
                12'd3875: logsin <= 24'd02065119;
                12'd3876: logsin <= 24'd02065405;
                12'd3877: logsin <= 24'd02065690;
                12'd3878: logsin <= 24'd02065974;
                12'd3879: logsin <= 24'd02066256;
                12'd3880: logsin <= 24'd02066538;
                12'd3881: logsin <= 24'd02066818;
                12'd3882: logsin <= 24'd02067096;
                12'd3883: logsin <= 24'd02067374;
                12'd3884: logsin <= 24'd02067650;
                12'd3885: logsin <= 24'd02067925;
                12'd3886: logsin <= 24'd02068199;
                12'd3887: logsin <= 24'd02068472;
                12'd3888: logsin <= 24'd02068743;
                12'd3889: logsin <= 24'd02069013;
                12'd3890: logsin <= 24'd02069282;
                12'd3891: logsin <= 24'd02069549;
                12'd3892: logsin <= 24'd02069816;
                12'd3893: logsin <= 24'd02070081;
                12'd3894: logsin <= 24'd02070345;
                12'd3895: logsin <= 24'd02070607;
                12'd3896: logsin <= 24'd02070869;
                12'd3897: logsin <= 24'd02071129;
                12'd3898: logsin <= 24'd02071387;
                12'd3899: logsin <= 24'd02071645;
                12'd3900: logsin <= 24'd02071901;
                12'd3901: logsin <= 24'd02072156;
                12'd3902: logsin <= 24'd02072410;
                12'd3903: logsin <= 24'd02072663;
                12'd3904: logsin <= 24'd02072914;
                12'd3905: logsin <= 24'd02073164;
                12'd3906: logsin <= 24'd02073413;
                12'd3907: logsin <= 24'd02073660;
                12'd3908: logsin <= 24'd02073907;
                12'd3909: logsin <= 24'd02074152;
                12'd3910: logsin <= 24'd02074395;
                12'd3911: logsin <= 24'd02074638;
                12'd3912: logsin <= 24'd02074879;
                12'd3913: logsin <= 24'd02075119;
                12'd3914: logsin <= 24'd02075358;
                12'd3915: logsin <= 24'd02075595;
                12'd3916: logsin <= 24'd02075831;
                12'd3917: logsin <= 24'd02076066;
                12'd3918: logsin <= 24'd02076300;
                12'd3919: logsin <= 24'd02076532;
                12'd3920: logsin <= 24'd02076763;
                12'd3921: logsin <= 24'd02076993;
                12'd3922: logsin <= 24'd02077222;
                12'd3923: logsin <= 24'd02077449;
                12'd3924: logsin <= 24'd02077675;
                12'd3925: logsin <= 24'd02077900;
                12'd3926: logsin <= 24'd02078123;
                12'd3927: logsin <= 24'd02078345;
                12'd3928: logsin <= 24'd02078566;
                12'd3929: logsin <= 24'd02078786;
                12'd3930: logsin <= 24'd02079004;
                12'd3931: logsin <= 24'd02079221;
                12'd3932: logsin <= 24'd02079437;
                12'd3933: logsin <= 24'd02079651;
                12'd3934: logsin <= 24'd02079865;
                12'd3935: logsin <= 24'd02080077;
                12'd3936: logsin <= 24'd02080287;
                12'd3937: logsin <= 24'd02080497;
                12'd3938: logsin <= 24'd02080705;
                12'd3939: logsin <= 24'd02080912;
                12'd3940: logsin <= 24'd02081117;
                12'd3941: logsin <= 24'd02081321;
                12'd3942: logsin <= 24'd02081524;
                12'd3943: logsin <= 24'd02081726;
                12'd3944: logsin <= 24'd02081926;
                12'd3945: logsin <= 24'd02082125;
                12'd3946: logsin <= 24'd02082323;
                12'd3947: logsin <= 24'd02082520;
                12'd3948: logsin <= 24'd02082715;
                12'd3949: logsin <= 24'd02082909;
                12'd3950: logsin <= 24'd02083102;
                12'd3951: logsin <= 24'd02083293;
                12'd3952: logsin <= 24'd02083483;
                12'd3953: logsin <= 24'd02083672;
                12'd3954: logsin <= 24'd02083860;
                12'd3955: logsin <= 24'd02084046;
                12'd3956: logsin <= 24'd02084231;
                12'd3957: logsin <= 24'd02084414;
                12'd3958: logsin <= 24'd02084597;
                12'd3959: logsin <= 24'd02084778;
                12'd3960: logsin <= 24'd02084957;
                12'd3961: logsin <= 24'd02085136;
                12'd3962: logsin <= 24'd02085313;
                12'd3963: logsin <= 24'd02085489;
                12'd3964: logsin <= 24'd02085664;
                12'd3965: logsin <= 24'd02085837;
                12'd3966: logsin <= 24'd02086009;
                12'd3967: logsin <= 24'd02086179;
                12'd3968: logsin <= 24'd02086349;
                12'd3969: logsin <= 24'd02086517;
                12'd3970: logsin <= 24'd02086684;
                12'd3971: logsin <= 24'd02086849;
                12'd3972: logsin <= 24'd02087013;
                12'd3973: logsin <= 24'd02087176;
                12'd3974: logsin <= 24'd02087338;
                12'd3975: logsin <= 24'd02087498;
                12'd3976: logsin <= 24'd02087657;
                12'd3977: logsin <= 24'd02087815;
                12'd3978: logsin <= 24'd02087971;
                12'd3979: logsin <= 24'd02088126;
                12'd3980: logsin <= 24'd02088280;
                12'd3981: logsin <= 24'd02088432;
                12'd3982: logsin <= 24'd02088583;
                12'd3983: logsin <= 24'd02088733;
                12'd3984: logsin <= 24'd02088881;
                12'd3985: logsin <= 24'd02089029;
                12'd3986: logsin <= 24'd02089175;
                12'd3987: logsin <= 24'd02089319;
                12'd3988: logsin <= 24'd02089462;
                12'd3989: logsin <= 24'd02089604;
                12'd3990: logsin <= 24'd02089745;
                12'd3991: logsin <= 24'd02089884;
                12'd3992: logsin <= 24'd02090022;
                12'd3993: logsin <= 24'd02090159;
                12'd3994: logsin <= 24'd02090294;
                12'd3995: logsin <= 24'd02090429;
                12'd3996: logsin <= 24'd02090561;
                12'd3997: logsin <= 24'd02090693;
                12'd3998: logsin <= 24'd02090823;
                12'd3999: logsin <= 24'd02090952;
                12'd4000: logsin <= 24'd02091079;
                12'd4001: logsin <= 24'd02091205;
                12'd4002: logsin <= 24'd02091330;
                12'd4003: logsin <= 24'd02091454;
                12'd4004: logsin <= 24'd02091576;
                12'd4005: logsin <= 24'd02091697;
                12'd4006: logsin <= 24'd02091817;
                12'd4007: logsin <= 24'd02091935;
                12'd4008: logsin <= 24'd02092052;
                12'd4009: logsin <= 24'd02092168;
                12'd4010: logsin <= 24'd02092282;
                12'd4011: logsin <= 24'd02092395;
                12'd4012: logsin <= 24'd02092507;
                12'd4013: logsin <= 24'd02092617;
                12'd4014: logsin <= 24'd02092726;
                12'd4015: logsin <= 24'd02092834;
                12'd4016: logsin <= 24'd02092940;
                12'd4017: logsin <= 24'd02093045;
                12'd4018: logsin <= 24'd02093149;
                12'd4019: logsin <= 24'd02093252;
                12'd4020: logsin <= 24'd02093353;
                12'd4021: logsin <= 24'd02093453;
                12'd4022: logsin <= 24'd02093551;
                12'd4023: logsin <= 24'd02093648;
                12'd4024: logsin <= 24'd02093744;
                12'd4025: logsin <= 24'd02093839;
                12'd4026: logsin <= 24'd02093932;
                12'd4027: logsin <= 24'd02094024;
                12'd4028: logsin <= 24'd02094114;
                12'd4029: logsin <= 24'd02094204;
                12'd4030: logsin <= 24'd02094291;
                12'd4031: logsin <= 24'd02094378;
                12'd4032: logsin <= 24'd02094463;
                12'd4033: logsin <= 24'd02094547;
                12'd4034: logsin <= 24'd02094630;
                12'd4035: logsin <= 24'd02094711;
                12'd4036: logsin <= 24'd02094791;
                12'd4037: logsin <= 24'd02094870;
                12'd4038: logsin <= 24'd02094947;
                12'd4039: logsin <= 24'd02095023;
                12'd4040: logsin <= 24'd02095097;
                12'd4041: logsin <= 24'd02095171;
                12'd4042: logsin <= 24'd02095243;
                12'd4043: logsin <= 24'd02095313;
                12'd4044: logsin <= 24'd02095383;
                12'd4045: logsin <= 24'd02095451;
                12'd4046: logsin <= 24'd02095517;
                12'd4047: logsin <= 24'd02095583;
                12'd4048: logsin <= 24'd02095647;
                12'd4049: logsin <= 24'd02095709;
                12'd4050: logsin <= 24'd02095771;
                12'd4051: logsin <= 24'd02095831;
                12'd4052: logsin <= 24'd02095889;
                12'd4053: logsin <= 24'd02095947;
                12'd4054: logsin <= 24'd02096003;
                12'd4055: logsin <= 24'd02096057;
                12'd4056: logsin <= 24'd02096111;
                12'd4057: logsin <= 24'd02096163;
                12'd4058: logsin <= 24'd02096213;
                12'd4059: logsin <= 24'd02096263;
                12'd4060: logsin <= 24'd02096311;
                12'd4061: logsin <= 24'd02096357;
                12'd4062: logsin <= 24'd02096403;
                12'd4063: logsin <= 24'd02096447;
                12'd4064: logsin <= 24'd02096490;
                12'd4065: logsin <= 24'd02096531;
                12'd4066: logsin <= 24'd02096571;
                12'd4067: logsin <= 24'd02096610;
                12'd4068: logsin <= 24'd02096647;
                12'd4069: logsin <= 24'd02096683;
                12'd4070: logsin <= 24'd02096718;
                12'd4071: logsin <= 24'd02096751;
                12'd4072: logsin <= 24'd02096783;
                12'd4073: logsin <= 24'd02096814;
                12'd4074: logsin <= 24'd02096843;
                12'd4075: logsin <= 24'd02096871;
                12'd4076: logsin <= 24'd02096898;
                12'd4077: logsin <= 24'd02096923;
                12'd4078: logsin <= 24'd02096947;
                12'd4079: logsin <= 24'd02096970;
                12'd4080: logsin <= 24'd02096991;
                12'd4081: logsin <= 24'd02097011;
                12'd4082: logsin <= 24'd02097030;
                12'd4083: logsin <= 24'd02097047;
                12'd4084: logsin <= 24'd02097063;
                12'd4085: logsin <= 24'd02097078;
                12'd4086: logsin <= 24'd02097091;
                12'd4087: logsin <= 24'd02097103;
                12'd4088: logsin <= 24'd02097114;
                12'd4089: logsin <= 24'd02097123;
                12'd4090: logsin <= 24'd02097131;
                12'd4091: logsin <= 24'd02097138;
                12'd4092: logsin <= 24'd02097143;
                12'd4093: logsin <= 24'd02097147;
                12'd4094: logsin <= 24'd02097150;
                12'd4095: logsin <= 24'd02097151;
            endcase
        4'b10: //clean512 12/24-bit
            case (addr[15:4])
                12'd0000: logsin <= 24'd00000000;
                12'd0001: logsin <= 24'd00000000;
                12'd0002: logsin <= 24'd00000001;
                12'd0003: logsin <= 24'd00000003;
                12'd0004: logsin <= 24'd00000005;
                12'd0005: logsin <= 24'd00000008;
                12'd0006: logsin <= 24'd00000011;
                12'd0007: logsin <= 24'd00000015;
                12'd0008: logsin <= 24'd00000020;
                12'd0009: logsin <= 24'd00000025;
                12'd0010: logsin <= 24'd00000031;
                12'd0011: logsin <= 24'd00000037;
                12'd0012: logsin <= 24'd00000044;
                12'd0013: logsin <= 24'd00000052;
                12'd0014: logsin <= 24'd00000060;
                12'd0015: logsin <= 24'd00000069;
                12'd0016: logsin <= 24'd00000079;
                12'd0017: logsin <= 24'd00000089;
                12'd0018: logsin <= 24'd00000100;
                12'd0019: logsin <= 24'd00000111;
                12'd0020: logsin <= 24'd00000123;
                12'd0021: logsin <= 24'd00000136;
                12'd0022: logsin <= 24'd00000149;
                12'd0023: logsin <= 24'd00000163;
                12'd0024: logsin <= 24'd00000178;
                12'd0025: logsin <= 24'd00000193;
                12'd0026: logsin <= 24'd00000208;
                12'd0027: logsin <= 24'd00000225;
                12'd0028: logsin <= 24'd00000242;
                12'd0029: logsin <= 24'd00000259;
                12'd0030: logsin <= 24'd00000278;
                12'd0031: logsin <= 24'd00000296;
                12'd0032: logsin <= 24'd00000316;
                12'd0033: logsin <= 24'd00000336;
                12'd0034: logsin <= 24'd00000357;
                12'd0035: logsin <= 24'd00000378;
                12'd0036: logsin <= 24'd00000400;
                12'd0037: logsin <= 24'd00000422;
                12'd0038: logsin <= 24'd00000445;
                12'd0039: logsin <= 24'd00000469;
                12'd0040: logsin <= 24'd00000493;
                12'd0041: logsin <= 24'd00000518;
                12'd0042: logsin <= 24'd00000544;
                12'd0043: logsin <= 24'd00000570;
                12'd0044: logsin <= 24'd00000597;
                12'd0045: logsin <= 24'd00000624;
                12'd0046: logsin <= 24'd00000653;
                12'd0047: logsin <= 24'd00000681;
                12'd0048: logsin <= 24'd00000711;
                12'd0049: logsin <= 24'd00000740;
                12'd0050: logsin <= 24'd00000771;
                12'd0051: logsin <= 24'd00000802;
                12'd0052: logsin <= 24'd00000834;
                12'd0053: logsin <= 24'd00000866;
                12'd0054: logsin <= 24'd00000899;
                12'd0055: logsin <= 24'd00000933;
                12'd0056: logsin <= 24'd00000967;
                12'd0057: logsin <= 24'd00001002;
                12'd0058: logsin <= 24'd00001037;
                12'd0059: logsin <= 24'd00001073;
                12'd0060: logsin <= 24'd00001110;
                12'd0061: logsin <= 24'd00001147;
                12'd0062: logsin <= 24'd00001185;
                12'd0063: logsin <= 24'd00001224;
                12'd0064: logsin <= 24'd00001263;
                12'd0065: logsin <= 24'd00001303;
                12'd0066: logsin <= 24'd00001343;
                12'd0067: logsin <= 24'd00001384;
                12'd0068: logsin <= 24'd00001426;
                12'd0069: logsin <= 24'd00001468;
                12'd0070: logsin <= 24'd00001511;
                12'd0071: logsin <= 24'd00001554;
                12'd0072: logsin <= 24'd00001598;
                12'd0073: logsin <= 24'd00001643;
                12'd0074: logsin <= 24'd00001688;
                12'd0075: logsin <= 24'd00001734;
                12'd0076: logsin <= 24'd00001781;
                12'd0077: logsin <= 24'd00001828;
                12'd0078: logsin <= 24'd00001876;
                12'd0079: logsin <= 24'd00001924;
                12'd0080: logsin <= 24'd00001973;
                12'd0081: logsin <= 24'd00002023;
                12'd0082: logsin <= 24'd00002073;
                12'd0083: logsin <= 24'd00002124;
                12'd0084: logsin <= 24'd00002175;
                12'd0085: logsin <= 24'd00002228;
                12'd0086: logsin <= 24'd00002280;
                12'd0087: logsin <= 24'd00002334;
                12'd0088: logsin <= 24'd00002388;
                12'd0089: logsin <= 24'd00002442;
                12'd0090: logsin <= 24'd00002497;
                12'd0091: logsin <= 24'd00002553;
                12'd0092: logsin <= 24'd00002609;
                12'd0093: logsin <= 24'd00002666;
                12'd0094: logsin <= 24'd00002724;
                12'd0095: logsin <= 24'd00002782;
                12'd0096: logsin <= 24'd00002841;
                12'd0097: logsin <= 24'd00002901;
                12'd0098: logsin <= 24'd00002961;
                12'd0099: logsin <= 24'd00003021;
                12'd0100: logsin <= 24'd00003083;
                12'd0101: logsin <= 24'd00003145;
                12'd0102: logsin <= 24'd00003207;
                12'd0103: logsin <= 24'd00003270;
                12'd0104: logsin <= 24'd00003334;
                12'd0105: logsin <= 24'd00003399;
                12'd0106: logsin <= 24'd00003464;
                12'd0107: logsin <= 24'd00003529;
                12'd0108: logsin <= 24'd00003595;
                12'd0109: logsin <= 24'd00003662;
                12'd0110: logsin <= 24'd00003730;
                12'd0111: logsin <= 24'd00003798;
                12'd0112: logsin <= 24'd00003867;
                12'd0113: logsin <= 24'd00003936;
                12'd0114: logsin <= 24'd00004006;
                12'd0115: logsin <= 24'd00004076;
                12'd0116: logsin <= 24'd00004147;
                12'd0117: logsin <= 24'd00004219;
                12'd0118: logsin <= 24'd00004292;
                12'd0119: logsin <= 24'd00004365;
                12'd0120: logsin <= 24'd00004438;
                12'd0121: logsin <= 24'd00004512;
                12'd0122: logsin <= 24'd00004587;
                12'd0123: logsin <= 24'd00004663;
                12'd0124: logsin <= 24'd00004739;
                12'd0125: logsin <= 24'd00004815;
                12'd0126: logsin <= 24'd00004893;
                12'd0127: logsin <= 24'd00004971;
                12'd0128: logsin <= 24'd00005049;
                12'd0129: logsin <= 24'd00005128;
                12'd0130: logsin <= 24'd00005208;
                12'd0131: logsin <= 24'd00005288;
                12'd0132: logsin <= 24'd00005369;
                12'd0133: logsin <= 24'd00005451;
                12'd0134: logsin <= 24'd00005533;
                12'd0135: logsin <= 24'd00005616;
                12'd0136: logsin <= 24'd00005699;
                12'd0137: logsin <= 24'd00005784;
                12'd0138: logsin <= 24'd00005868;
                12'd0139: logsin <= 24'd00005953;
                12'd0140: logsin <= 24'd00006039;
                12'd0141: logsin <= 24'd00006126;
                12'd0142: logsin <= 24'd00006213;
                12'd0143: logsin <= 24'd00006301;
                12'd0144: logsin <= 24'd00006389;
                12'd0145: logsin <= 24'd00006478;
                12'd0146: logsin <= 24'd00006568;
                12'd0147: logsin <= 24'd00006658;
                12'd0148: logsin <= 24'd00006748;
                12'd0149: logsin <= 24'd00006840;
                12'd0150: logsin <= 24'd00006932;
                12'd0151: logsin <= 24'd00007025;
                12'd0152: logsin <= 24'd00007118;
                12'd0153: logsin <= 24'd00007212;
                12'd0154: logsin <= 24'd00007306;
                12'd0155: logsin <= 24'd00007401;
                12'd0156: logsin <= 24'd00007497;
                12'd0157: logsin <= 24'd00007593;
                12'd0158: logsin <= 24'd00007690;
                12'd0159: logsin <= 24'd00007788;
                12'd0160: logsin <= 24'd00007886;
                12'd0161: logsin <= 24'd00007985;
                12'd0162: logsin <= 24'd00008084;
                12'd0163: logsin <= 24'd00008184;
                12'd0164: logsin <= 24'd00008284;
                12'd0165: logsin <= 24'd00008386;
                12'd0166: logsin <= 24'd00008487;
                12'd0167: logsin <= 24'd00008590;
                12'd0168: logsin <= 24'd00008693;
                12'd0169: logsin <= 24'd00008797;
                12'd0170: logsin <= 24'd00008901;
                12'd0171: logsin <= 24'd00009006;
                12'd0172: logsin <= 24'd00009111;
                12'd0173: logsin <= 24'd00009217;
                12'd0174: logsin <= 24'd00009324;
                12'd0175: logsin <= 24'd00009431;
                12'd0176: logsin <= 24'd00009539;
                12'd0177: logsin <= 24'd00009648;
                12'd0178: logsin <= 24'd00009757;
                12'd0179: logsin <= 24'd00009867;
                12'd0180: logsin <= 24'd00009977;
                12'd0181: logsin <= 24'd00010088;
                12'd0182: logsin <= 24'd00010200;
                12'd0183: logsin <= 24'd00010312;
                12'd0184: logsin <= 24'd00010425;
                12'd0185: logsin <= 24'd00010538;
                12'd0186: logsin <= 24'd00010652;
                12'd0187: logsin <= 24'd00010767;
                12'd0188: logsin <= 24'd00010882;
                12'd0189: logsin <= 24'd00010998;
                12'd0190: logsin <= 24'd00011114;
                12'd0191: logsin <= 24'd00011232;
                12'd0192: logsin <= 24'd00011349;
                12'd0193: logsin <= 24'd00011468;
                12'd0194: logsin <= 24'd00011586;
                12'd0195: logsin <= 24'd00011706;
                12'd0196: logsin <= 24'd00011826;
                12'd0197: logsin <= 24'd00011947;
                12'd0198: logsin <= 24'd00012068;
                12'd0199: logsin <= 24'd00012190;
                12'd0200: logsin <= 24'd00012313;
                12'd0201: logsin <= 24'd00012436;
                12'd0202: logsin <= 24'd00012560;
                12'd0203: logsin <= 24'd00012684;
                12'd0204: logsin <= 24'd00012809;
                12'd0205: logsin <= 24'd00012935;
                12'd0206: logsin <= 24'd00013061;
                12'd0207: logsin <= 24'd00013188;
                12'd0208: logsin <= 24'd00013315;
                12'd0209: logsin <= 24'd00013443;
                12'd0210: logsin <= 24'd00013572;
                12'd0211: logsin <= 24'd00013701;
                12'd0212: logsin <= 24'd00013831;
                12'd0213: logsin <= 24'd00013962;
                12'd0214: logsin <= 24'd00014093;
                12'd0215: logsin <= 24'd00014225;
                12'd0216: logsin <= 24'd00014357;
                12'd0217: logsin <= 24'd00014490;
                12'd0218: logsin <= 24'd00014623;
                12'd0219: logsin <= 24'd00014758;
                12'd0220: logsin <= 24'd00014892;
                12'd0221: logsin <= 24'd00015028;
                12'd0222: logsin <= 24'd00015164;
                12'd0223: logsin <= 24'd00015300;
                12'd0224: logsin <= 24'd00015438;
                12'd0225: logsin <= 24'd00015575;
                12'd0226: logsin <= 24'd00015714;
                12'd0227: logsin <= 24'd00015853;
                12'd0228: logsin <= 24'd00015992;
                12'd0229: logsin <= 24'd00016133;
                12'd0230: logsin <= 24'd00016273;
                12'd0231: logsin <= 24'd00016415;
                12'd0232: logsin <= 24'd00016557;
                12'd0233: logsin <= 24'd00016700;
                12'd0234: logsin <= 24'd00016843;
                12'd0235: logsin <= 24'd00016987;
                12'd0236: logsin <= 24'd00017131;
                12'd0237: logsin <= 24'd00017276;
                12'd0238: logsin <= 24'd00017422;
                12'd0239: logsin <= 24'd00017568;
                12'd0240: logsin <= 24'd00017715;
                12'd0241: logsin <= 24'd00017863;
                12'd0242: logsin <= 24'd00018011;
                12'd0243: logsin <= 24'd00018160;
                12'd0244: logsin <= 24'd00018309;
                12'd0245: logsin <= 24'd00018459;
                12'd0246: logsin <= 24'd00018609;
                12'd0247: logsin <= 24'd00018760;
                12'd0248: logsin <= 24'd00018912;
                12'd0249: logsin <= 24'd00019065;
                12'd0250: logsin <= 24'd00019218;
                12'd0251: logsin <= 24'd00019371;
                12'd0252: logsin <= 24'd00019525;
                12'd0253: logsin <= 24'd00019680;
                12'd0254: logsin <= 24'd00019836;
                12'd0255: logsin <= 24'd00019991;
                12'd0256: logsin <= 24'd00020148;
                12'd0257: logsin <= 24'd00020305;
                12'd0258: logsin <= 24'd00020463;
                12'd0259: logsin <= 24'd00020622;
                12'd0260: logsin <= 24'd00020781;
                12'd0261: logsin <= 24'd00020940;
                12'd0262: logsin <= 24'd00021100;
                12'd0263: logsin <= 24'd00021261;
                12'd0264: logsin <= 24'd00021423;
                12'd0265: logsin <= 24'd00021585;
                12'd0266: logsin <= 24'd00021747;
                12'd0267: logsin <= 24'd00021911;
                12'd0268: logsin <= 24'd00022074;
                12'd0269: logsin <= 24'd00022239;
                12'd0270: logsin <= 24'd00022404;
                12'd0271: logsin <= 24'd00022570;
                12'd0272: logsin <= 24'd00022736;
                12'd0273: logsin <= 24'd00022903;
                12'd0274: logsin <= 24'd00023070;
                12'd0275: logsin <= 24'd00023238;
                12'd0276: logsin <= 24'd00023407;
                12'd0277: logsin <= 24'd00023576;
                12'd0278: logsin <= 24'd00023746;
                12'd0279: logsin <= 24'd00023917;
                12'd0280: logsin <= 24'd00024088;
                12'd0281: logsin <= 24'd00024259;
                12'd0282: logsin <= 24'd00024432;
                12'd0283: logsin <= 24'd00024605;
                12'd0284: logsin <= 24'd00024778;
                12'd0285: logsin <= 24'd00024952;
                12'd0286: logsin <= 24'd00025127;
                12'd0287: logsin <= 24'd00025302;
                12'd0288: logsin <= 24'd00025478;
                12'd0289: logsin <= 24'd00025655;
                12'd0290: logsin <= 24'd00025832;
                12'd0291: logsin <= 24'd00026010;
                12'd0292: logsin <= 24'd00026188;
                12'd0293: logsin <= 24'd00026367;
                12'd0294: logsin <= 24'd00026546;
                12'd0295: logsin <= 24'd00026726;
                12'd0296: logsin <= 24'd00026907;
                12'd0297: logsin <= 24'd00027088;
                12'd0298: logsin <= 24'd00027270;
                12'd0299: logsin <= 24'd00027453;
                12'd0300: logsin <= 24'd00027636;
                12'd0301: logsin <= 24'd00027820;
                12'd0302: logsin <= 24'd00028004;
                12'd0303: logsin <= 24'd00028189;
                12'd0304: logsin <= 24'd00028375;
                12'd0305: logsin <= 24'd00028561;
                12'd0306: logsin <= 24'd00028747;
                12'd0307: logsin <= 24'd00028935;
                12'd0308: logsin <= 24'd00029123;
                12'd0309: logsin <= 24'd00029311;
                12'd0310: logsin <= 24'd00029500;
                12'd0311: logsin <= 24'd00029690;
                12'd0312: logsin <= 24'd00029880;
                12'd0313: logsin <= 24'd00030071;
                12'd0314: logsin <= 24'd00030263;
                12'd0315: logsin <= 24'd00030455;
                12'd0316: logsin <= 24'd00030648;
                12'd0317: logsin <= 24'd00030841;
                12'd0318: logsin <= 24'd00031035;
                12'd0319: logsin <= 24'd00031229;
                12'd0320: logsin <= 24'd00031425;
                12'd0321: logsin <= 24'd00031620;
                12'd0322: logsin <= 24'd00031817;
                12'd0323: logsin <= 24'd00032013;
                12'd0324: logsin <= 24'd00032211;
                12'd0325: logsin <= 24'd00032409;
                12'd0326: logsin <= 24'd00032608;
                12'd0327: logsin <= 24'd00032807;
                12'd0328: logsin <= 24'd00033007;
                12'd0329: logsin <= 24'd00033207;
                12'd0330: logsin <= 24'd00033409;
                12'd0331: logsin <= 24'd00033610;
                12'd0332: logsin <= 24'd00033813;
                12'd0333: logsin <= 24'd00034015;
                12'd0334: logsin <= 24'd00034219;
                12'd0335: logsin <= 24'd00034423;
                12'd0336: logsin <= 24'd00034628;
                12'd0337: logsin <= 24'd00034833;
                12'd0338: logsin <= 24'd00035039;
                12'd0339: logsin <= 24'd00035245;
                12'd0340: logsin <= 24'd00035452;
                12'd0341: logsin <= 24'd00035660;
                12'd0342: logsin <= 24'd00035868;
                12'd0343: logsin <= 24'd00036077;
                12'd0344: logsin <= 24'd00036287;
                12'd0345: logsin <= 24'd00036497;
                12'd0346: logsin <= 24'd00036707;
                12'd0347: logsin <= 24'd00036918;
                12'd0348: logsin <= 24'd00037130;
                12'd0349: logsin <= 24'd00037343;
                12'd0350: logsin <= 24'd00037556;
                12'd0351: logsin <= 24'd00037769;
                12'd0352: logsin <= 24'd00037984;
                12'd0353: logsin <= 24'd00038198;
                12'd0354: logsin <= 24'd00038414;
                12'd0355: logsin <= 24'd00038630;
                12'd0356: logsin <= 24'd00038846;
                12'd0357: logsin <= 24'd00039063;
                12'd0358: logsin <= 24'd00039281;
                12'd0359: logsin <= 24'd00039500;
                12'd0360: logsin <= 24'd00039719;
                12'd0361: logsin <= 24'd00039938;
                12'd0362: logsin <= 24'd00040158;
                12'd0363: logsin <= 24'd00040379;
                12'd0364: logsin <= 24'd00040600;
                12'd0365: logsin <= 24'd00040822;
                12'd0366: logsin <= 24'd00041045;
                12'd0367: logsin <= 24'd00041268;
                12'd0368: logsin <= 24'd00041492;
                12'd0369: logsin <= 24'd00041716;
                12'd0370: logsin <= 24'd00041941;
                12'd0371: logsin <= 24'd00042166;
                12'd0372: logsin <= 24'd00042392;
                12'd0373: logsin <= 24'd00042619;
                12'd0374: logsin <= 24'd00042846;
                12'd0375: logsin <= 24'd00043074;
                12'd0376: logsin <= 24'd00043303;
                12'd0377: logsin <= 24'd00043532;
                12'd0378: logsin <= 24'd00043761;
                12'd0379: logsin <= 24'd00043991;
                12'd0380: logsin <= 24'd00044222;
                12'd0381: logsin <= 24'd00044454;
                12'd0382: logsin <= 24'd00044686;
                12'd0383: logsin <= 24'd00044918;
                12'd0384: logsin <= 24'd00045151;
                12'd0385: logsin <= 24'd00045385;
                12'd0386: logsin <= 24'd00045619;
                12'd0387: logsin <= 24'd00045854;
                12'd0388: logsin <= 24'd00046090;
                12'd0389: logsin <= 24'd00046326;
                12'd0390: logsin <= 24'd00046563;
                12'd0391: logsin <= 24'd00046800;
                12'd0392: logsin <= 24'd00047038;
                12'd0393: logsin <= 24'd00047276;
                12'd0394: logsin <= 24'd00047515;
                12'd0395: logsin <= 24'd00047755;
                12'd0396: logsin <= 24'd00047995;
                12'd0397: logsin <= 24'd00048236;
                12'd0398: logsin <= 24'd00048478;
                12'd0399: logsin <= 24'd00048720;
                12'd0400: logsin <= 24'd00048962;
                12'd0401: logsin <= 24'd00049205;
                12'd0402: logsin <= 24'd00049449;
                12'd0403: logsin <= 24'd00049693;
                12'd0404: logsin <= 24'd00049938;
                12'd0405: logsin <= 24'd00050184;
                12'd0406: logsin <= 24'd00050430;
                12'd0407: logsin <= 24'd00050677;
                12'd0408: logsin <= 24'd00050924;
                12'd0409: logsin <= 24'd00051172;
                12'd0410: logsin <= 24'd00051420;
                12'd0411: logsin <= 24'd00051669;
                12'd0412: logsin <= 24'd00051919;
                12'd0413: logsin <= 24'd00052169;
                12'd0414: logsin <= 24'd00052420;
                12'd0415: logsin <= 24'd00052672;
                12'd0416: logsin <= 24'd00052924;
                12'd0417: logsin <= 24'd00053176;
                12'd0418: logsin <= 24'd00053429;
                12'd0419: logsin <= 24'd00053683;
                12'd0420: logsin <= 24'd00053937;
                12'd0421: logsin <= 24'd00054192;
                12'd0422: logsin <= 24'd00054448;
                12'd0423: logsin <= 24'd00054704;
                12'd0424: logsin <= 24'd00054960;
                12'd0425: logsin <= 24'd00055218;
                12'd0426: logsin <= 24'd00055476;
                12'd0427: logsin <= 24'd00055734;
                12'd0428: logsin <= 24'd00055993;
                12'd0429: logsin <= 24'd00056253;
                12'd0430: logsin <= 24'd00056513;
                12'd0431: logsin <= 24'd00056774;
                12'd0432: logsin <= 24'd00057035;
                12'd0433: logsin <= 24'd00057297;
                12'd0434: logsin <= 24'd00057559;
                12'd0435: logsin <= 24'd00057822;
                12'd0436: logsin <= 24'd00058086;
                12'd0437: logsin <= 24'd00058350;
                12'd0438: logsin <= 24'd00058615;
                12'd0439: logsin <= 24'd00058881;
                12'd0440: logsin <= 24'd00059147;
                12'd0441: logsin <= 24'd00059413;
                12'd0442: logsin <= 24'd00059680;
                12'd0443: logsin <= 24'd00059948;
                12'd0444: logsin <= 24'd00060216;
                12'd0445: logsin <= 24'd00060485;
                12'd0446: logsin <= 24'd00060755;
                12'd0447: logsin <= 24'd00061025;
                12'd0448: logsin <= 24'd00061295;
                12'd0449: logsin <= 24'd00061567;
                12'd0450: logsin <= 24'd00061839;
                12'd0451: logsin <= 24'd00062111;
                12'd0452: logsin <= 24'd00062384;
                12'd0453: logsin <= 24'd00062657;
                12'd0454: logsin <= 24'd00062932;
                12'd0455: logsin <= 24'd00063206;
                12'd0456: logsin <= 24'd00063482;
                12'd0457: logsin <= 24'd00063757;
                12'd0458: logsin <= 24'd00064034;
                12'd0459: logsin <= 24'd00064311;
                12'd0460: logsin <= 24'd00064589;
                12'd0461: logsin <= 24'd00064867;
                12'd0462: logsin <= 24'd00065146;
                12'd0463: logsin <= 24'd00065425;
                12'd0464: logsin <= 24'd00065705;
                12'd0465: logsin <= 24'd00065985;
                12'd0466: logsin <= 24'd00066266;
                12'd0467: logsin <= 24'd00066548;
                12'd0468: logsin <= 24'd00066830;
                12'd0469: logsin <= 24'd00067113;
                12'd0470: logsin <= 24'd00067396;
                12'd0471: logsin <= 24'd00067680;
                12'd0472: logsin <= 24'd00067965;
                12'd0473: logsin <= 24'd00068250;
                12'd0474: logsin <= 24'd00068536;
                12'd0475: logsin <= 24'd00068822;
                12'd0476: logsin <= 24'd00069109;
                12'd0477: logsin <= 24'd00069396;
                12'd0478: logsin <= 24'd00069684;
                12'd0479: logsin <= 24'd00069973;
                12'd0480: logsin <= 24'd00070262;
                12'd0481: logsin <= 24'd00070552;
                12'd0482: logsin <= 24'd00070842;
                12'd0483: logsin <= 24'd00071133;
                12'd0484: logsin <= 24'd00071425;
                12'd0485: logsin <= 24'd00071717;
                12'd0486: logsin <= 24'd00072009;
                12'd0487: logsin <= 24'd00072302;
                12'd0488: logsin <= 24'd00072596;
                12'd0489: logsin <= 24'd00072890;
                12'd0490: logsin <= 24'd00073185;
                12'd0491: logsin <= 24'd00073481;
                12'd0492: logsin <= 24'd00073777;
                12'd0493: logsin <= 24'd00074073;
                12'd0494: logsin <= 24'd00074371;
                12'd0495: logsin <= 24'd00074668;
                12'd0496: logsin <= 24'd00074967;
                12'd0497: logsin <= 24'd00075266;
                12'd0498: logsin <= 24'd00075565;
                12'd0499: logsin <= 24'd00075865;
                12'd0500: logsin <= 24'd00076166;
                12'd0501: logsin <= 24'd00076467;
                12'd0502: logsin <= 24'd00076769;
                12'd0503: logsin <= 24'd00077071;
                12'd0504: logsin <= 24'd00077374;
                12'd0505: logsin <= 24'd00077678;
                12'd0506: logsin <= 24'd00077982;
                12'd0507: logsin <= 24'd00078286;
                12'd0508: logsin <= 24'd00078592;
                12'd0509: logsin <= 24'd00078897;
                12'd0510: logsin <= 24'd00079204;
                12'd0511: logsin <= 24'd00079511;
                12'd0512: logsin <= 24'd00079818;
                12'd0513: logsin <= 24'd00080126;
                12'd0514: logsin <= 24'd00080435;
                12'd0515: logsin <= 24'd00080744;
                12'd0516: logsin <= 24'd00081054;
                12'd0517: logsin <= 24'd00081364;
                12'd0518: logsin <= 24'd00081675;
                12'd0519: logsin <= 24'd00081986;
                12'd0520: logsin <= 24'd00082298;
                12'd0521: logsin <= 24'd00082611;
                12'd0522: logsin <= 24'd00082924;
                12'd0523: logsin <= 24'd00083238;
                12'd0524: logsin <= 24'd00083552;
                12'd0525: logsin <= 24'd00083867;
                12'd0526: logsin <= 24'd00084183;
                12'd0527: logsin <= 24'd00084499;
                12'd0528: logsin <= 24'd00084815;
                12'd0529: logsin <= 24'd00085132;
                12'd0530: logsin <= 24'd00085450;
                12'd0531: logsin <= 24'd00085768;
                12'd0532: logsin <= 24'd00086087;
                12'd0533: logsin <= 24'd00086407;
                12'd0534: logsin <= 24'd00086727;
                12'd0535: logsin <= 24'd00087047;
                12'd0536: logsin <= 24'd00087368;
                12'd0537: logsin <= 24'd00087690;
                12'd0538: logsin <= 24'd00088012;
                12'd0539: logsin <= 24'd00088335;
                12'd0540: logsin <= 24'd00088658;
                12'd0541: logsin <= 24'd00088982;
                12'd0542: logsin <= 24'd00089307;
                12'd0543: logsin <= 24'd00089632;
                12'd0544: logsin <= 24'd00089958;
                12'd0545: logsin <= 24'd00090284;
                12'd0546: logsin <= 24'd00090611;
                12'd0547: logsin <= 24'd00090938;
                12'd0548: logsin <= 24'd00091266;
                12'd0549: logsin <= 24'd00091594;
                12'd0550: logsin <= 24'd00091923;
                12'd0551: logsin <= 24'd00092253;
                12'd0552: logsin <= 24'd00092583;
                12'd0553: logsin <= 24'd00092914;
                12'd0554: logsin <= 24'd00093245;
                12'd0555: logsin <= 24'd00093577;
                12'd0556: logsin <= 24'd00093909;
                12'd0557: logsin <= 24'd00094242;
                12'd0558: logsin <= 24'd00094576;
                12'd0559: logsin <= 24'd00094910;
                12'd0560: logsin <= 24'd00095244;
                12'd0561: logsin <= 24'd00095579;
                12'd0562: logsin <= 24'd00095915;
                12'd0563: logsin <= 24'd00096252;
                12'd0564: logsin <= 24'd00096588;
                12'd0565: logsin <= 24'd00096926;
                12'd0566: logsin <= 24'd00097264;
                12'd0567: logsin <= 24'd00097602;
                12'd0568: logsin <= 24'd00097942;
                12'd0569: logsin <= 24'd00098281;
                12'd0570: logsin <= 24'd00098621;
                12'd0571: logsin <= 24'd00098962;
                12'd0572: logsin <= 24'd00099304;
                12'd0573: logsin <= 24'd00099645;
                12'd0574: logsin <= 24'd00099988;
                12'd0575: logsin <= 24'd00100331;
                12'd0576: logsin <= 24'd00100675;
                12'd0577: logsin <= 24'd00101019;
                12'd0578: logsin <= 24'd00101363;
                12'd0579: logsin <= 24'd00101709;
                12'd0580: logsin <= 24'd00102054;
                12'd0581: logsin <= 24'd00102401;
                12'd0582: logsin <= 24'd00102748;
                12'd0583: logsin <= 24'd00103095;
                12'd0584: logsin <= 24'd00103443;
                12'd0585: logsin <= 24'd00103792;
                12'd0586: logsin <= 24'd00104141;
                12'd0587: logsin <= 24'd00104491;
                12'd0588: logsin <= 24'd00104841;
                12'd0589: logsin <= 24'd00105192;
                12'd0590: logsin <= 24'd00105543;
                12'd0591: logsin <= 24'd00105895;
                12'd0592: logsin <= 24'd00106248;
                12'd0593: logsin <= 24'd00106601;
                12'd0594: logsin <= 24'd00106954;
                12'd0595: logsin <= 24'd00107308;
                12'd0596: logsin <= 24'd00107663;
                12'd0597: logsin <= 24'd00108018;
                12'd0598: logsin <= 24'd00108374;
                12'd0599: logsin <= 24'd00108730;
                12'd0600: logsin <= 24'd00109087;
                12'd0601: logsin <= 24'd00109445;
                12'd0602: logsin <= 24'd00109803;
                12'd0603: logsin <= 24'd00110161;
                12'd0604: logsin <= 24'd00110520;
                12'd0605: logsin <= 24'd00110880;
                12'd0606: logsin <= 24'd00111240;
                12'd0607: logsin <= 24'd00111601;
                12'd0608: logsin <= 24'd00111962;
                12'd0609: logsin <= 24'd00112324;
                12'd0610: logsin <= 24'd00112687;
                12'd0611: logsin <= 24'd00113050;
                12'd0612: logsin <= 24'd00113413;
                12'd0613: logsin <= 24'd00113777;
                12'd0614: logsin <= 24'd00114142;
                12'd0615: logsin <= 24'd00114507;
                12'd0616: logsin <= 24'd00114873;
                12'd0617: logsin <= 24'd00115239;
                12'd0618: logsin <= 24'd00115606;
                12'd0619: logsin <= 24'd00115973;
                12'd0620: logsin <= 24'd00116341;
                12'd0621: logsin <= 24'd00116710;
                12'd0622: logsin <= 24'd00117079;
                12'd0623: logsin <= 24'd00117448;
                12'd0624: logsin <= 24'd00117818;
                12'd0625: logsin <= 24'd00118189;
                12'd0626: logsin <= 24'd00118560;
                12'd0627: logsin <= 24'd00118932;
                12'd0628: logsin <= 24'd00119304;
                12'd0629: logsin <= 24'd00119677;
                12'd0630: logsin <= 24'd00120051;
                12'd0631: logsin <= 24'd00120425;
                12'd0632: logsin <= 24'd00120799;
                12'd0633: logsin <= 24'd00121174;
                12'd0634: logsin <= 24'd00121550;
                12'd0635: logsin <= 24'd00121926;
                12'd0636: logsin <= 24'd00122302;
                12'd0637: logsin <= 24'd00122680;
                12'd0638: logsin <= 24'd00123057;
                12'd0639: logsin <= 24'd00123436;
                12'd0640: logsin <= 24'd00123815;
                12'd0641: logsin <= 24'd00124194;
                12'd0642: logsin <= 24'd00124574;
                12'd0643: logsin <= 24'd00124954;
                12'd0644: logsin <= 24'd00125335;
                12'd0645: logsin <= 24'd00125717;
                12'd0646: logsin <= 24'd00126099;
                12'd0647: logsin <= 24'd00126482;
                12'd0648: logsin <= 24'd00126865;
                12'd0649: logsin <= 24'd00127249;
                12'd0650: logsin <= 24'd00127633;
                12'd0651: logsin <= 24'd00128018;
                12'd0652: logsin <= 24'd00128403;
                12'd0653: logsin <= 24'd00128789;
                12'd0654: logsin <= 24'd00129175;
                12'd0655: logsin <= 24'd00129562;
                12'd0656: logsin <= 24'd00129950;
                12'd0657: logsin <= 24'd00130338;
                12'd0658: logsin <= 24'd00130727;
                12'd0659: logsin <= 24'd00131116;
                12'd0660: logsin <= 24'd00131505;
                12'd0661: logsin <= 24'd00131896;
                12'd0662: logsin <= 24'd00132286;
                12'd0663: logsin <= 24'd00132678;
                12'd0664: logsin <= 24'd00133070;
                12'd0665: logsin <= 24'd00133462;
                12'd0666: logsin <= 24'd00133855;
                12'd0667: logsin <= 24'd00134248;
                12'd0668: logsin <= 24'd00134642;
                12'd0669: logsin <= 24'd00135037;
                12'd0670: logsin <= 24'd00135432;
                12'd0671: logsin <= 24'd00135828;
                12'd0672: logsin <= 24'd00136224;
                12'd0673: logsin <= 24'd00136620;
                12'd0674: logsin <= 24'd00137018;
                12'd0675: logsin <= 24'd00137415;
                12'd0676: logsin <= 24'd00137814;
                12'd0677: logsin <= 24'd00138212;
                12'd0678: logsin <= 24'd00138612;
                12'd0679: logsin <= 24'd00139012;
                12'd0680: logsin <= 24'd00139412;
                12'd0681: logsin <= 24'd00139813;
                12'd0682: logsin <= 24'd00140215;
                12'd0683: logsin <= 24'd00140617;
                12'd0684: logsin <= 24'd00141019;
                12'd0685: logsin <= 24'd00141422;
                12'd0686: logsin <= 24'd00141826;
                12'd0687: logsin <= 24'd00142230;
                12'd0688: logsin <= 24'd00142635;
                12'd0689: logsin <= 24'd00143040;
                12'd0690: logsin <= 24'd00143446;
                12'd0691: logsin <= 24'd00143852;
                12'd0692: logsin <= 24'd00144259;
                12'd0693: logsin <= 24'd00144666;
                12'd0694: logsin <= 24'd00145074;
                12'd0695: logsin <= 24'd00145483;
                12'd0696: logsin <= 24'd00145892;
                12'd0697: logsin <= 24'd00146301;
                12'd0698: logsin <= 24'd00146711;
                12'd0699: logsin <= 24'd00147122;
                12'd0700: logsin <= 24'd00147533;
                12'd0701: logsin <= 24'd00147944;
                12'd0702: logsin <= 24'd00148356;
                12'd0703: logsin <= 24'd00148769;
                12'd0704: logsin <= 24'd00149182;
                12'd0705: logsin <= 24'd00149596;
                12'd0706: logsin <= 24'd00150010;
                12'd0707: logsin <= 24'd00150425;
                12'd0708: logsin <= 24'd00150840;
                12'd0709: logsin <= 24'd00151256;
                12'd0710: logsin <= 24'd00151673;
                12'd0711: logsin <= 24'd00152090;
                12'd0712: logsin <= 24'd00152507;
                12'd0713: logsin <= 24'd00152925;
                12'd0714: logsin <= 24'd00153343;
                12'd0715: logsin <= 24'd00153762;
                12'd0716: logsin <= 24'd00154182;
                12'd0717: logsin <= 24'd00154602;
                12'd0718: logsin <= 24'd00155023;
                12'd0719: logsin <= 24'd00155444;
                12'd0720: logsin <= 24'd00155865;
                12'd0721: logsin <= 24'd00156288;
                12'd0722: logsin <= 24'd00156710;
                12'd0723: logsin <= 24'd00157133;
                12'd0724: logsin <= 24'd00157557;
                12'd0725: logsin <= 24'd00157981;
                12'd0726: logsin <= 24'd00158406;
                12'd0727: logsin <= 24'd00158832;
                12'd0728: logsin <= 24'd00159257;
                12'd0729: logsin <= 24'd00159684;
                12'd0730: logsin <= 24'd00160111;
                12'd0731: logsin <= 24'd00160538;
                12'd0732: logsin <= 24'd00160966;
                12'd0733: logsin <= 24'd00161394;
                12'd0734: logsin <= 24'd00161823;
                12'd0735: logsin <= 24'd00162253;
                12'd0736: logsin <= 24'd00162683;
                12'd0737: logsin <= 24'd00163113;
                12'd0738: logsin <= 24'd00163544;
                12'd0739: logsin <= 24'd00163976;
                12'd0740: logsin <= 24'd00164408;
                12'd0741: logsin <= 24'd00164841;
                12'd0742: logsin <= 24'd00165274;
                12'd0743: logsin <= 24'd00165707;
                12'd0744: logsin <= 24'd00166142;
                12'd0745: logsin <= 24'd00166576;
                12'd0746: logsin <= 24'd00167012;
                12'd0747: logsin <= 24'd00167447;
                12'd0748: logsin <= 24'd00167884;
                12'd0749: logsin <= 24'd00168320;
                12'd0750: logsin <= 24'd00168758;
                12'd0751: logsin <= 24'd00169195;
                12'd0752: logsin <= 24'd00169634;
                12'd0753: logsin <= 24'd00170073;
                12'd0754: logsin <= 24'd00170512;
                12'd0755: logsin <= 24'd00170952;
                12'd0756: logsin <= 24'd00171392;
                12'd0757: logsin <= 24'd00171833;
                12'd0758: logsin <= 24'd00172274;
                12'd0759: logsin <= 24'd00172716;
                12'd0760: logsin <= 24'd00173159;
                12'd0761: logsin <= 24'd00173602;
                12'd0762: logsin <= 24'd00174045;
                12'd0763: logsin <= 24'd00174489;
                12'd0764: logsin <= 24'd00174934;
                12'd0765: logsin <= 24'd00175379;
                12'd0766: logsin <= 24'd00175824;
                12'd0767: logsin <= 24'd00176270;
                12'd0768: logsin <= 24'd00176717;
                12'd0769: logsin <= 24'd00177164;
                12'd0770: logsin <= 24'd00177612;
                12'd0771: logsin <= 24'd00178060;
                12'd0772: logsin <= 24'd00178508;
                12'd0773: logsin <= 24'd00178957;
                12'd0774: logsin <= 24'd00179407;
                12'd0775: logsin <= 24'd00179857;
                12'd0776: logsin <= 24'd00180308;
                12'd0777: logsin <= 24'd00180759;
                12'd0778: logsin <= 24'd00181211;
                12'd0779: logsin <= 24'd00181663;
                12'd0780: logsin <= 24'd00182116;
                12'd0781: logsin <= 24'd00182569;
                12'd0782: logsin <= 24'd00183022;
                12'd0783: logsin <= 24'd00183477;
                12'd0784: logsin <= 24'd00183931;
                12'd0785: logsin <= 24'd00184387;
                12'd0786: logsin <= 24'd00184842;
                12'd0787: logsin <= 24'd00185299;
                12'd0788: logsin <= 24'd00185755;
                12'd0789: logsin <= 24'd00186213;
                12'd0790: logsin <= 24'd00186671;
                12'd0791: logsin <= 24'd00187129;
                12'd0792: logsin <= 24'd00187588;
                12'd0793: logsin <= 24'd00188047;
                12'd0794: logsin <= 24'd00188507;
                12'd0795: logsin <= 24'd00188967;
                12'd0796: logsin <= 24'd00189428;
                12'd0797: logsin <= 24'd00189889;
                12'd0798: logsin <= 24'd00190351;
                12'd0799: logsin <= 24'd00190813;
                12'd0800: logsin <= 24'd00191276;
                12'd0801: logsin <= 24'd00191740;
                12'd0802: logsin <= 24'd00192203;
                12'd0803: logsin <= 24'd00192668;
                12'd0804: logsin <= 24'd00193133;
                12'd0805: logsin <= 24'd00193598;
                12'd0806: logsin <= 24'd00194064;
                12'd0807: logsin <= 24'd00194530;
                12'd0808: logsin <= 24'd00194997;
                12'd0809: logsin <= 24'd00195464;
                12'd0810: logsin <= 24'd00195932;
                12'd0811: logsin <= 24'd00196401;
                12'd0812: logsin <= 24'd00196870;
                12'd0813: logsin <= 24'd00197339;
                12'd0814: logsin <= 24'd00197809;
                12'd0815: logsin <= 24'd00198279;
                12'd0816: logsin <= 24'd00198750;
                12'd0817: logsin <= 24'd00199221;
                12'd0818: logsin <= 24'd00199693;
                12'd0819: logsin <= 24'd00200166;
                12'd0820: logsin <= 24'd00200639;
                12'd0821: logsin <= 24'd00201112;
                12'd0822: logsin <= 24'd00201586;
                12'd0823: logsin <= 24'd00202060;
                12'd0824: logsin <= 24'd00202535;
                12'd0825: logsin <= 24'd00203010;
                12'd0826: logsin <= 24'd00203486;
                12'd0827: logsin <= 24'd00203963;
                12'd0828: logsin <= 24'd00204439;
                12'd0829: logsin <= 24'd00204917;
                12'd0830: logsin <= 24'd00205395;
                12'd0831: logsin <= 24'd00205873;
                12'd0832: logsin <= 24'd00206352;
                12'd0833: logsin <= 24'd00206831;
                12'd0834: logsin <= 24'd00207311;
                12'd0835: logsin <= 24'd00207791;
                12'd0836: logsin <= 24'd00208272;
                12'd0837: logsin <= 24'd00208753;
                12'd0838: logsin <= 24'd00209235;
                12'd0839: logsin <= 24'd00209718;
                12'd0840: logsin <= 24'd00210200;
                12'd0841: logsin <= 24'd00210684;
                12'd0842: logsin <= 24'd00211167;
                12'd0843: logsin <= 24'd00211652;
                12'd0844: logsin <= 24'd00212137;
                12'd0845: logsin <= 24'd00212622;
                12'd0846: logsin <= 24'd00213108;
                12'd0847: logsin <= 24'd00213594;
                12'd0848: logsin <= 24'd00214081;
                12'd0849: logsin <= 24'd00214568;
                12'd0850: logsin <= 24'd00215055;
                12'd0851: logsin <= 24'd00215544;
                12'd0852: logsin <= 24'd00216032;
                12'd0853: logsin <= 24'd00216522;
                12'd0854: logsin <= 24'd00217011;
                12'd0855: logsin <= 24'd00217501;
                12'd0856: logsin <= 24'd00217992;
                12'd0857: logsin <= 24'd00218483;
                12'd0858: logsin <= 24'd00218975;
                12'd0859: logsin <= 24'd00219467;
                12'd0860: logsin <= 24'd00219960;
                12'd0861: logsin <= 24'd00220453;
                12'd0862: logsin <= 24'd00220946;
                12'd0863: logsin <= 24'd00221440;
                12'd0864: logsin <= 24'd00221935;
                12'd0865: logsin <= 24'd00222430;
                12'd0866: logsin <= 24'd00222925;
                12'd0867: logsin <= 24'd00223421;
                12'd0868: logsin <= 24'd00223918;
                12'd0869: logsin <= 24'd00224415;
                12'd0870: logsin <= 24'd00224912;
                12'd0871: logsin <= 24'd00225410;
                12'd0872: logsin <= 24'd00225909;
                12'd0873: logsin <= 24'd00226408;
                12'd0874: logsin <= 24'd00226907;
                12'd0875: logsin <= 24'd00227407;
                12'd0876: logsin <= 24'd00227907;
                12'd0877: logsin <= 24'd00228408;
                12'd0878: logsin <= 24'd00228910;
                12'd0879: logsin <= 24'd00229411;
                12'd0880: logsin <= 24'd00229914;
                12'd0881: logsin <= 24'd00230416;
                12'd0882: logsin <= 24'd00230920;
                12'd0883: logsin <= 24'd00231423;
                12'd0884: logsin <= 24'd00231928;
                12'd0885: logsin <= 24'd00232432;
                12'd0886: logsin <= 24'd00232938;
                12'd0887: logsin <= 24'd00233443;
                12'd0888: logsin <= 24'd00233949;
                12'd0889: logsin <= 24'd00234456;
                12'd0890: logsin <= 24'd00234963;
                12'd0891: logsin <= 24'd00235471;
                12'd0892: logsin <= 24'd00235979;
                12'd0893: logsin <= 24'd00236487;
                12'd0894: logsin <= 24'd00236996;
                12'd0895: logsin <= 24'd00237506;
                12'd0896: logsin <= 24'd00238016;
                12'd0897: logsin <= 24'd00238526;
                12'd0898: logsin <= 24'd00239037;
                12'd0899: logsin <= 24'd00239549;
                12'd0900: logsin <= 24'd00240060;
                12'd0901: logsin <= 24'd00240573;
                12'd0902: logsin <= 24'd00241086;
                12'd0903: logsin <= 24'd00241599;
                12'd0904: logsin <= 24'd00242113;
                12'd0905: logsin <= 24'd00242627;
                12'd0906: logsin <= 24'd00243142;
                12'd0907: logsin <= 24'd00243657;
                12'd0908: logsin <= 24'd00244173;
                12'd0909: logsin <= 24'd00244689;
                12'd0910: logsin <= 24'd00245205;
                12'd0911: logsin <= 24'd00245722;
                12'd0912: logsin <= 24'd00246240;
                12'd0913: logsin <= 24'd00246758;
                12'd0914: logsin <= 24'd00247277;
                12'd0915: logsin <= 24'd00247795;
                12'd0916: logsin <= 24'd00248315;
                12'd0917: logsin <= 24'd00248835;
                12'd0918: logsin <= 24'd00249355;
                12'd0919: logsin <= 24'd00249876;
                12'd0920: logsin <= 24'd00250397;
                12'd0921: logsin <= 24'd00250919;
                12'd0922: logsin <= 24'd00251442;
                12'd0923: logsin <= 24'd00251964;
                12'd0924: logsin <= 24'd00252487;
                12'd0925: logsin <= 24'd00253011;
                12'd0926: logsin <= 24'd00253535;
                12'd0927: logsin <= 24'd00254060;
                12'd0928: logsin <= 24'd00254585;
                12'd0929: logsin <= 24'd00255111;
                12'd0930: logsin <= 24'd00255637;
                12'd0931: logsin <= 24'd00256163;
                12'd0932: logsin <= 24'd00256690;
                12'd0933: logsin <= 24'd00257217;
                12'd0934: logsin <= 24'd00257745;
                12'd0935: logsin <= 24'd00258274;
                12'd0936: logsin <= 24'd00258802;
                12'd0937: logsin <= 24'd00259332;
                12'd0938: logsin <= 24'd00259861;
                12'd0939: logsin <= 24'd00260392;
                12'd0940: logsin <= 24'd00260922;
                12'd0941: logsin <= 24'd00261453;
                12'd0942: logsin <= 24'd00261985;
                12'd0943: logsin <= 24'd00262517;
                12'd0944: logsin <= 24'd00263050;
                12'd0945: logsin <= 24'd00263583;
                12'd0946: logsin <= 24'd00264116;
                12'd0947: logsin <= 24'd00264650;
                12'd0948: logsin <= 24'd00265184;
                12'd0949: logsin <= 24'd00265719;
                12'd0950: logsin <= 24'd00266254;
                12'd0951: logsin <= 24'd00266790;
                12'd0952: logsin <= 24'd00267326;
                12'd0953: logsin <= 24'd00267863;
                12'd0954: logsin <= 24'd00268400;
                12'd0955: logsin <= 24'd00268938;
                12'd0956: logsin <= 24'd00269476;
                12'd0957: logsin <= 24'd00270014;
                12'd0958: logsin <= 24'd00270553;
                12'd0959: logsin <= 24'd00271093;
                12'd0960: logsin <= 24'd00271632;
                12'd0961: logsin <= 24'd00272173;
                12'd0962: logsin <= 24'd00272714;
                12'd0963: logsin <= 24'd00273255;
                12'd0964: logsin <= 24'd00273796;
                12'd0965: logsin <= 24'd00274339;
                12'd0966: logsin <= 24'd00274881;
                12'd0967: logsin <= 24'd00275424;
                12'd0968: logsin <= 24'd00275968;
                12'd0969: logsin <= 24'd00276512;
                12'd0970: logsin <= 24'd00277056;
                12'd0971: logsin <= 24'd00277601;
                12'd0972: logsin <= 24'd00278146;
                12'd0973: logsin <= 24'd00278692;
                12'd0974: logsin <= 24'd00279238;
                12'd0975: logsin <= 24'd00279785;
                12'd0976: logsin <= 24'd00280332;
                12'd0977: logsin <= 24'd00280880;
                12'd0978: logsin <= 24'd00281428;
                12'd0979: logsin <= 24'd00281976;
                12'd0980: logsin <= 24'd00282525;
                12'd0981: logsin <= 24'd00283075;
                12'd0982: logsin <= 24'd00283625;
                12'd0983: logsin <= 24'd00284175;
                12'd0984: logsin <= 24'd00284726;
                12'd0985: logsin <= 24'd00285277;
                12'd0986: logsin <= 24'd00285829;
                12'd0987: logsin <= 24'd00286381;
                12'd0988: logsin <= 24'd00286933;
                12'd0989: logsin <= 24'd00287486;
                12'd0990: logsin <= 24'd00288040;
                12'd0991: logsin <= 24'd00288594;
                12'd0992: logsin <= 24'd00289148;
                12'd0993: logsin <= 24'd00289703;
                12'd0994: logsin <= 24'd00290258;
                12'd0995: logsin <= 24'd00290814;
                12'd0996: logsin <= 24'd00291370;
                12'd0997: logsin <= 24'd00291926;
                12'd0998: logsin <= 24'd00292483;
                12'd0999: logsin <= 24'd00293041;
                12'd1000: logsin <= 24'd00293599;
                12'd1001: logsin <= 24'd00294157;
                12'd1002: logsin <= 24'd00294716;
                12'd1003: logsin <= 24'd00295275;
                12'd1004: logsin <= 24'd00295835;
                12'd1005: logsin <= 24'd00296395;
                12'd1006: logsin <= 24'd00296955;
                12'd1007: logsin <= 24'd00297516;
                12'd1008: logsin <= 24'd00298078;
                12'd1009: logsin <= 24'd00298640;
                12'd1010: logsin <= 24'd00299202;
                12'd1011: logsin <= 24'd00299765;
                12'd1012: logsin <= 24'd00300328;
                12'd1013: logsin <= 24'd00300892;
                12'd1014: logsin <= 24'd00301456;
                12'd1015: logsin <= 24'd00302020;
                12'd1016: logsin <= 24'd00302585;
                12'd1017: logsin <= 24'd00303151;
                12'd1018: logsin <= 24'd00303717;
                12'd1019: logsin <= 24'd00304283;
                12'd1020: logsin <= 24'd00304850;
                12'd1021: logsin <= 24'd00305417;
                12'd1022: logsin <= 24'd00305984;
                12'd1023: logsin <= 24'd00306552;
                12'd1024: logsin <= 24'd00307121;
                12'd1025: logsin <= 24'd00307690;
                12'd1026: logsin <= 24'd00308259;
                12'd1027: logsin <= 24'd00308829;
                12'd1028: logsin <= 24'd00309399;
                12'd1029: logsin <= 24'd00309970;
                12'd1030: logsin <= 24'd00310541;
                12'd1031: logsin <= 24'd00311112;
                12'd1032: logsin <= 24'd00311684;
                12'd1033: logsin <= 24'd00312257;
                12'd1034: logsin <= 24'd00312829;
                12'd1035: logsin <= 24'd00313403;
                12'd1036: logsin <= 24'd00313976;
                12'd1037: logsin <= 24'd00314550;
                12'd1038: logsin <= 24'd00315125;
                12'd1039: logsin <= 24'd00315700;
                12'd1040: logsin <= 24'd00316275;
                12'd1041: logsin <= 24'd00316851;
                12'd1042: logsin <= 24'd00317428;
                12'd1043: logsin <= 24'd00318004;
                12'd1044: logsin <= 24'd00318581;
                12'd1045: logsin <= 24'd00319159;
                12'd1046: logsin <= 24'd00319737;
                12'd1047: logsin <= 24'd00320315;
                12'd1048: logsin <= 24'd00320894;
                12'd1049: logsin <= 24'd00321473;
                12'd1050: logsin <= 24'd00322053;
                12'd1051: logsin <= 24'd00322633;
                12'd1052: logsin <= 24'd00323214;
                12'd1053: logsin <= 24'd00323795;
                12'd1054: logsin <= 24'd00324376;
                12'd1055: logsin <= 24'd00324958;
                12'd1056: logsin <= 24'd00325540;
                12'd1057: logsin <= 24'd00326123;
                12'd1058: logsin <= 24'd00326706;
                12'd1059: logsin <= 24'd00327290;
                12'd1060: logsin <= 24'd00327874;
                12'd1061: logsin <= 24'd00328458;
                12'd1062: logsin <= 24'd00329043;
                12'd1063: logsin <= 24'd00329628;
                12'd1064: logsin <= 24'd00330214;
                12'd1065: logsin <= 24'd00330800;
                12'd1066: logsin <= 24'd00331386;
                12'd1067: logsin <= 24'd00331973;
                12'd1068: logsin <= 24'd00332561;
                12'd1069: logsin <= 24'd00333148;
                12'd1070: logsin <= 24'd00333736;
                12'd1071: logsin <= 24'd00334325;
                12'd1072: logsin <= 24'd00334914;
                12'd1073: logsin <= 24'd00335504;
                12'd1074: logsin <= 24'd00336093;
                12'd1075: logsin <= 24'd00336684;
                12'd1076: logsin <= 24'd00337274;
                12'd1077: logsin <= 24'd00337866;
                12'd1078: logsin <= 24'd00338457;
                12'd1079: logsin <= 24'd00339049;
                12'd1080: logsin <= 24'd00339641;
                12'd1081: logsin <= 24'd00340234;
                12'd1082: logsin <= 24'd00340827;
                12'd1083: logsin <= 24'd00341421;
                12'd1084: logsin <= 24'd00342015;
                12'd1085: logsin <= 24'd00342610;
                12'd1086: logsin <= 24'd00343204;
                12'd1087: logsin <= 24'd00343800;
                12'd1088: logsin <= 24'd00344395;
                12'd1089: logsin <= 24'd00344992;
                12'd1090: logsin <= 24'd00345588;
                12'd1091: logsin <= 24'd00346185;
                12'd1092: logsin <= 24'd00346782;
                12'd1093: logsin <= 24'd00347380;
                12'd1094: logsin <= 24'd00347978;
                12'd1095: logsin <= 24'd00348577;
                12'd1096: logsin <= 24'd00349176;
                12'd1097: logsin <= 24'd00349775;
                12'd1098: logsin <= 24'd00350375;
                12'd1099: logsin <= 24'd00350975;
                12'd1100: logsin <= 24'd00351576;
                12'd1101: logsin <= 24'd00352177;
                12'd1102: logsin <= 24'd00352779;
                12'd1103: logsin <= 24'd00353380;
                12'd1104: logsin <= 24'd00353983;
                12'd1105: logsin <= 24'd00354585;
                12'd1106: logsin <= 24'd00355189;
                12'd1107: logsin <= 24'd00355792;
                12'd1108: logsin <= 24'd00356396;
                12'd1109: logsin <= 24'd00357000;
                12'd1110: logsin <= 24'd00357605;
                12'd1111: logsin <= 24'd00358210;
                12'd1112: logsin <= 24'd00358816;
                12'd1113: logsin <= 24'd00359422;
                12'd1114: logsin <= 24'd00360028;
                12'd1115: logsin <= 24'd00360635;
                12'd1116: logsin <= 24'd00361242;
                12'd1117: logsin <= 24'd00361849;
                12'd1118: logsin <= 24'd00362457;
                12'd1119: logsin <= 24'd00363066;
                12'd1120: logsin <= 24'd00363675;
                12'd1121: logsin <= 24'd00364284;
                12'd1122: logsin <= 24'd00364893;
                12'd1123: logsin <= 24'd00365503;
                12'd1124: logsin <= 24'd00366114;
                12'd1125: logsin <= 24'd00366725;
                12'd1126: logsin <= 24'd00367336;
                12'd1127: logsin <= 24'd00367947;
                12'd1128: logsin <= 24'd00368559;
                12'd1129: logsin <= 24'd00369172;
                12'd1130: logsin <= 24'd00369785;
                12'd1131: logsin <= 24'd00370398;
                12'd1132: logsin <= 24'd00371011;
                12'd1133: logsin <= 24'd00371625;
                12'd1134: logsin <= 24'd00372240;
                12'd1135: logsin <= 24'd00372855;
                12'd1136: logsin <= 24'd00373470;
                12'd1137: logsin <= 24'd00374085;
                12'd1138: logsin <= 24'd00374701;
                12'd1139: logsin <= 24'd00375318;
                12'd1140: logsin <= 24'd00375934;
                12'd1141: logsin <= 24'd00376552;
                12'd1142: logsin <= 24'd00377169;
                12'd1143: logsin <= 24'd00377787;
                12'd1144: logsin <= 24'd00378405;
                12'd1145: logsin <= 24'd00379024;
                12'd1146: logsin <= 24'd00379643;
                12'd1147: logsin <= 24'd00380263;
                12'd1148: logsin <= 24'd00380883;
                12'd1149: logsin <= 24'd00381503;
                12'd1150: logsin <= 24'd00382124;
                12'd1151: logsin <= 24'd00382745;
                12'd1152: logsin <= 24'd00383366;
                12'd1153: logsin <= 24'd00383988;
                12'd1154: logsin <= 24'd00384611;
                12'd1155: logsin <= 24'd00385233;
                12'd1156: logsin <= 24'd00385856;
                12'd1157: logsin <= 24'd00386480;
                12'd1158: logsin <= 24'd00387104;
                12'd1159: logsin <= 24'd00387728;
                12'd1160: logsin <= 24'd00388352;
                12'd1161: logsin <= 24'd00388977;
                12'd1162: logsin <= 24'd00389603;
                12'd1163: logsin <= 24'd00390229;
                12'd1164: logsin <= 24'd00390855;
                12'd1165: logsin <= 24'd00391481;
                12'd1166: logsin <= 24'd00392108;
                12'd1167: logsin <= 24'd00392736;
                12'd1168: logsin <= 24'd00393363;
                12'd1169: logsin <= 24'd00393991;
                12'd1170: logsin <= 24'd00394620;
                12'd1171: logsin <= 24'd00395249;
                12'd1172: logsin <= 24'd00395878;
                12'd1173: logsin <= 24'd00396508;
                12'd1174: logsin <= 24'd00397138;
                12'd1175: logsin <= 24'd00397768;
                12'd1176: logsin <= 24'd00398399;
                12'd1177: logsin <= 24'd00399030;
                12'd1178: logsin <= 24'd00399662;
                12'd1179: logsin <= 24'd00400294;
                12'd1180: logsin <= 24'd00400926;
                12'd1181: logsin <= 24'd00401559;
                12'd1182: logsin <= 24'd00402192;
                12'd1183: logsin <= 24'd00402825;
                12'd1184: logsin <= 24'd00403459;
                12'd1185: logsin <= 24'd00404093;
                12'd1186: logsin <= 24'd00404728;
                12'd1187: logsin <= 24'd00405363;
                12'd1188: logsin <= 24'd00405998;
                12'd1189: logsin <= 24'd00406634;
                12'd1190: logsin <= 24'd00407270;
                12'd1191: logsin <= 24'd00407906;
                12'd1192: logsin <= 24'd00408543;
                12'd1193: logsin <= 24'd00409180;
                12'd1194: logsin <= 24'd00409818;
                12'd1195: logsin <= 24'd00410456;
                12'd1196: logsin <= 24'd00411094;
                12'd1197: logsin <= 24'd00411733;
                12'd1198: logsin <= 24'd00412372;
                12'd1199: logsin <= 24'd00413012;
                12'd1200: logsin <= 24'd00413652;
                12'd1201: logsin <= 24'd00414292;
                12'd1202: logsin <= 24'd00414933;
                12'd1203: logsin <= 24'd00415573;
                12'd1204: logsin <= 24'd00416215;
                12'd1205: logsin <= 24'd00416857;
                12'd1206: logsin <= 24'd00417499;
                12'd1207: logsin <= 24'd00418141;
                12'd1208: logsin <= 24'd00418784;
                12'd1209: logsin <= 24'd00419427;
                12'd1210: logsin <= 24'd00420071;
                12'd1211: logsin <= 24'd00420715;
                12'd1212: logsin <= 24'd00421359;
                12'd1213: logsin <= 24'd00422004;
                12'd1214: logsin <= 24'd00422649;
                12'd1215: logsin <= 24'd00423294;
                12'd1216: logsin <= 24'd00423940;
                12'd1217: logsin <= 24'd00424586;
                12'd1218: logsin <= 24'd00425233;
                12'd1219: logsin <= 24'd00425880;
                12'd1220: logsin <= 24'd00426527;
                12'd1221: logsin <= 24'd00427174;
                12'd1222: logsin <= 24'd00427822;
                12'd1223: logsin <= 24'd00428471;
                12'd1224: logsin <= 24'd00429120;
                12'd1225: logsin <= 24'd00429769;
                12'd1226: logsin <= 24'd00430418;
                12'd1227: logsin <= 24'd00431068;
                12'd1228: logsin <= 24'd00431718;
                12'd1229: logsin <= 24'd00432369;
                12'd1230: logsin <= 24'd00433020;
                12'd1231: logsin <= 24'd00433671;
                12'd1232: logsin <= 24'd00434322;
                12'd1233: logsin <= 24'd00434974;
                12'd1234: logsin <= 24'd00435627;
                12'd1235: logsin <= 24'd00436279;
                12'd1236: logsin <= 24'd00436933;
                12'd1237: logsin <= 24'd00437586;
                12'd1238: logsin <= 24'd00438240;
                12'd1239: logsin <= 24'd00438894;
                12'd1240: logsin <= 24'd00439548;
                12'd1241: logsin <= 24'd00440203;
                12'd1242: logsin <= 24'd00440859;
                12'd1243: logsin <= 24'd00441514;
                12'd1244: logsin <= 24'd00442170;
                12'd1245: logsin <= 24'd00442826;
                12'd1246: logsin <= 24'd00443483;
                12'd1247: logsin <= 24'd00444140;
                12'd1248: logsin <= 24'd00444797;
                12'd1249: logsin <= 24'd00445455;
                12'd1250: logsin <= 24'd00446113;
                12'd1251: logsin <= 24'd00446772;
                12'd1252: logsin <= 24'd00447430;
                12'd1253: logsin <= 24'd00448089;
                12'd1254: logsin <= 24'd00448749;
                12'd1255: logsin <= 24'd00449409;
                12'd1256: logsin <= 24'd00450069;
                12'd1257: logsin <= 24'd00450730;
                12'd1258: logsin <= 24'd00451390;
                12'd1259: logsin <= 24'd00452052;
                12'd1260: logsin <= 24'd00452713;
                12'd1261: logsin <= 24'd00453375;
                12'd1262: logsin <= 24'd00454038;
                12'd1263: logsin <= 24'd00454700;
                12'd1264: logsin <= 24'd00455363;
                12'd1265: logsin <= 24'd00456027;
                12'd1266: logsin <= 24'd00456690;
                12'd1267: logsin <= 24'd00457354;
                12'd1268: logsin <= 24'd00458019;
                12'd1269: logsin <= 24'd00458683;
                12'd1270: logsin <= 24'd00459349;
                12'd1271: logsin <= 24'd00460014;
                12'd1272: logsin <= 24'd00460680;
                12'd1273: logsin <= 24'd00461346;
                12'd1274: logsin <= 24'd00462012;
                12'd1275: logsin <= 24'd00462679;
                12'd1276: logsin <= 24'd00463346;
                12'd1277: logsin <= 24'd00464014;
                12'd1278: logsin <= 24'd00464682;
                12'd1279: logsin <= 24'd00465350;
                12'd1280: logsin <= 24'd00466018;
                12'd1281: logsin <= 24'd00466687;
                12'd1282: logsin <= 24'd00467356;
                12'd1283: logsin <= 24'd00468026;
                12'd1284: logsin <= 24'd00468696;
                12'd1285: logsin <= 24'd00469366;
                12'd1286: logsin <= 24'd00470037;
                12'd1287: logsin <= 24'd00470708;
                12'd1288: logsin <= 24'd00471379;
                12'd1289: logsin <= 24'd00472051;
                12'd1290: logsin <= 24'd00472723;
                12'd1291: logsin <= 24'd00473395;
                12'd1292: logsin <= 24'd00474067;
                12'd1293: logsin <= 24'd00474740;
                12'd1294: logsin <= 24'd00475414;
                12'd1295: logsin <= 24'd00476087;
                12'd1296: logsin <= 24'd00476761;
                12'd1297: logsin <= 24'd00477436;
                12'd1298: logsin <= 24'd00478110;
                12'd1299: logsin <= 24'd00478785;
                12'd1300: logsin <= 24'd00479461;
                12'd1301: logsin <= 24'd00480136;
                12'd1302: logsin <= 24'd00480812;
                12'd1303: logsin <= 24'd00481489;
                12'd1304: logsin <= 24'd00482165;
                12'd1305: logsin <= 24'd00482842;
                12'd1306: logsin <= 24'd00483519;
                12'd1307: logsin <= 24'd00484197;
                12'd1308: logsin <= 24'd00484875;
                12'd1309: logsin <= 24'd00485553;
                12'd1310: logsin <= 24'd00486232;
                12'd1311: logsin <= 24'd00486911;
                12'd1312: logsin <= 24'd00487590;
                12'd1313: logsin <= 24'd00488270;
                12'd1314: logsin <= 24'd00488950;
                12'd1315: logsin <= 24'd00489630;
                12'd1316: logsin <= 24'd00490311;
                12'd1317: logsin <= 24'd00490992;
                12'd1318: logsin <= 24'd00491673;
                12'd1319: logsin <= 24'd00492355;
                12'd1320: logsin <= 24'd00493037;
                12'd1321: logsin <= 24'd00493719;
                12'd1322: logsin <= 24'd00494401;
                12'd1323: logsin <= 24'd00495084;
                12'd1324: logsin <= 24'd00495768;
                12'd1325: logsin <= 24'd00496451;
                12'd1326: logsin <= 24'd00497135;
                12'd1327: logsin <= 24'd00497819;
                12'd1328: logsin <= 24'd00498504;
                12'd1329: logsin <= 24'd00499189;
                12'd1330: logsin <= 24'd00499874;
                12'd1331: logsin <= 24'd00500559;
                12'd1332: logsin <= 24'd00501245;
                12'd1333: logsin <= 24'd00501931;
                12'd1334: logsin <= 24'd00502618;
                12'd1335: logsin <= 24'd00503305;
                12'd1336: logsin <= 24'd00503992;
                12'd1337: logsin <= 24'd00504679;
                12'd1338: logsin <= 24'd00505367;
                12'd1339: logsin <= 24'd00506055;
                12'd1340: logsin <= 24'd00506743;
                12'd1341: logsin <= 24'd00507432;
                12'd1342: logsin <= 24'd00508121;
                12'd1343: logsin <= 24'd00508811;
                12'd1344: logsin <= 24'd00509500;
                12'd1345: logsin <= 24'd00510190;
                12'd1346: logsin <= 24'd00510880;
                12'd1347: logsin <= 24'd00511571;
                12'd1348: logsin <= 24'd00512262;
                12'd1349: logsin <= 24'd00512953;
                12'd1350: logsin <= 24'd00513645;
                12'd1351: logsin <= 24'd00514337;
                12'd1352: logsin <= 24'd00515029;
                12'd1353: logsin <= 24'd00515721;
                12'd1354: logsin <= 24'd00516414;
                12'd1355: logsin <= 24'd00517107;
                12'd1356: logsin <= 24'd00517801;
                12'd1357: logsin <= 24'd00518495;
                12'd1358: logsin <= 24'd00519189;
                12'd1359: logsin <= 24'd00519883;
                12'd1360: logsin <= 24'd00520578;
                12'd1361: logsin <= 24'd00521273;
                12'd1362: logsin <= 24'd00521968;
                12'd1363: logsin <= 24'd00522664;
                12'd1364: logsin <= 24'd00523360;
                12'd1365: logsin <= 24'd00524056;
                12'd1366: logsin <= 24'd00524752;
                12'd1367: logsin <= 24'd00525449;
                12'd1368: logsin <= 24'd00526146;
                12'd1369: logsin <= 24'd00526844;
                12'd1370: logsin <= 24'd00527542;
                12'd1371: logsin <= 24'd00528240;
                12'd1372: logsin <= 24'd00528938;
                12'd1373: logsin <= 24'd00529637;
                12'd1374: logsin <= 24'd00530336;
                12'd1375: logsin <= 24'd00531035;
                12'd1376: logsin <= 24'd00531735;
                12'd1377: logsin <= 24'd00532435;
                12'd1378: logsin <= 24'd00533135;
                12'd1379: logsin <= 24'd00533835;
                12'd1380: logsin <= 24'd00534536;
                12'd1381: logsin <= 24'd00535237;
                12'd1382: logsin <= 24'd00535939;
                12'd1383: logsin <= 24'd00536641;
                12'd1384: logsin <= 24'd00537343;
                12'd1385: logsin <= 24'd00538045;
                12'd1386: logsin <= 24'd00538748;
                12'd1387: logsin <= 24'd00539451;
                12'd1388: logsin <= 24'd00540154;
                12'd1389: logsin <= 24'd00540857;
                12'd1390: logsin <= 24'd00541561;
                12'd1391: logsin <= 24'd00542265;
                12'd1392: logsin <= 24'd00542970;
                12'd1393: logsin <= 24'd00543674;
                12'd1394: logsin <= 24'd00544379;
                12'd1395: logsin <= 24'd00545085;
                12'd1396: logsin <= 24'd00545790;
                12'd1397: logsin <= 24'd00546496;
                12'd1398: logsin <= 24'd00547202;
                12'd1399: logsin <= 24'd00547909;
                12'd1400: logsin <= 24'd00548616;
                12'd1401: logsin <= 24'd00549323;
                12'd1402: logsin <= 24'd00550030;
                12'd1403: logsin <= 24'd00550738;
                12'd1404: logsin <= 24'd00551446;
                12'd1405: logsin <= 24'd00552154;
                12'd1406: logsin <= 24'd00552863;
                12'd1407: logsin <= 24'd00553572;
                12'd1408: logsin <= 24'd00554281;
                12'd1409: logsin <= 24'd00554990;
                12'd1410: logsin <= 24'd00555700;
                12'd1411: logsin <= 24'd00556410;
                12'd1412: logsin <= 24'd00557120;
                12'd1413: logsin <= 24'd00557831;
                12'd1414: logsin <= 24'd00558542;
                12'd1415: logsin <= 24'd00559253;
                12'd1416: logsin <= 24'd00559964;
                12'd1417: logsin <= 24'd00560676;
                12'd1418: logsin <= 24'd00561388;
                12'd1419: logsin <= 24'd00562100;
                12'd1420: logsin <= 24'd00562813;
                12'd1421: logsin <= 24'd00563526;
                12'd1422: logsin <= 24'd00564239;
                12'd1423: logsin <= 24'd00564952;
                12'd1424: logsin <= 24'd00565666;
                12'd1425: logsin <= 24'd00566380;
                12'd1426: logsin <= 24'd00567094;
                12'd1427: logsin <= 24'd00567809;
                12'd1428: logsin <= 24'd00568524;
                12'd1429: logsin <= 24'd00569239;
                12'd1430: logsin <= 24'd00569955;
                12'd1431: logsin <= 24'd00570670;
                12'd1432: logsin <= 24'd00571386;
                12'd1433: logsin <= 24'd00572103;
                12'd1434: logsin <= 24'd00572819;
                12'd1435: logsin <= 24'd00573536;
                12'd1436: logsin <= 24'd00574253;
                12'd1437: logsin <= 24'd00574970;
                12'd1438: logsin <= 24'd00575688;
                12'd1439: logsin <= 24'd00576406;
                12'd1440: logsin <= 24'd00577124;
                12'd1441: logsin <= 24'd00577843;
                12'd1442: logsin <= 24'd00578562;
                12'd1443: logsin <= 24'd00579281;
                12'd1444: logsin <= 24'd00580000;
                12'd1445: logsin <= 24'd00580720;
                12'd1446: logsin <= 24'd00581440;
                12'd1447: logsin <= 24'd00582160;
                12'd1448: logsin <= 24'd00582880;
                12'd1449: logsin <= 24'd00583601;
                12'd1450: logsin <= 24'd00584322;
                12'd1451: logsin <= 24'd00585043;
                12'd1452: logsin <= 24'd00585765;
                12'd1453: logsin <= 24'd00586486;
                12'd1454: logsin <= 24'd00587209;
                12'd1455: logsin <= 24'd00587931;
                12'd1456: logsin <= 24'd00588654;
                12'd1457: logsin <= 24'd00589376;
                12'd1458: logsin <= 24'd00590100;
                12'd1459: logsin <= 24'd00590823;
                12'd1460: logsin <= 24'd00591547;
                12'd1461: logsin <= 24'd00592271;
                12'd1462: logsin <= 24'd00592995;
                12'd1463: logsin <= 24'd00593719;
                12'd1464: logsin <= 24'd00594444;
                12'd1465: logsin <= 24'd00595169;
                12'd1466: logsin <= 24'd00595895;
                12'd1467: logsin <= 24'd00596620;
                12'd1468: logsin <= 24'd00597346;
                12'd1469: logsin <= 24'd00598072;
                12'd1470: logsin <= 24'd00598798;
                12'd1471: logsin <= 24'd00599525;
                12'd1472: logsin <= 24'd00600252;
                12'd1473: logsin <= 24'd00600979;
                12'd1474: logsin <= 24'd00601707;
                12'd1475: logsin <= 24'd00602434;
                12'd1476: logsin <= 24'd00603162;
                12'd1477: logsin <= 24'd00603890;
                12'd1478: logsin <= 24'd00604619;
                12'd1479: logsin <= 24'd00605348;
                12'd1480: logsin <= 24'd00606077;
                12'd1481: logsin <= 24'd00606806;
                12'd1482: logsin <= 24'd00607535;
                12'd1483: logsin <= 24'd00608265;
                12'd1484: logsin <= 24'd00608995;
                12'd1485: logsin <= 24'd00609726;
                12'd1486: logsin <= 24'd00610456;
                12'd1487: logsin <= 24'd00611187;
                12'd1488: logsin <= 24'd00611918;
                12'd1489: logsin <= 24'd00612649;
                12'd1490: logsin <= 24'd00613381;
                12'd1491: logsin <= 24'd00614113;
                12'd1492: logsin <= 24'd00614845;
                12'd1493: logsin <= 24'd00615577;
                12'd1494: logsin <= 24'd00616310;
                12'd1495: logsin <= 24'd00617043;
                12'd1496: logsin <= 24'd00617776;
                12'd1497: logsin <= 24'd00618509;
                12'd1498: logsin <= 24'd00619243;
                12'd1499: logsin <= 24'd00619977;
                12'd1500: logsin <= 24'd00620711;
                12'd1501: logsin <= 24'd00621445;
                12'd1502: logsin <= 24'd00622180;
                12'd1503: logsin <= 24'd00622915;
                12'd1504: logsin <= 24'd00623650;
                12'd1505: logsin <= 24'd00624385;
                12'd1506: logsin <= 24'd00625121;
                12'd1507: logsin <= 24'd00625857;
                12'd1508: logsin <= 24'd00626593;
                12'd1509: logsin <= 24'd00627329;
                12'd1510: logsin <= 24'd00628066;
                12'd1511: logsin <= 24'd00628803;
                12'd1512: logsin <= 24'd00629540;
                12'd1513: logsin <= 24'd00630277;
                12'd1514: logsin <= 24'd00631015;
                12'd1515: logsin <= 24'd00631752;
                12'd1516: logsin <= 24'd00632491;
                12'd1517: logsin <= 24'd00633229;
                12'd1518: logsin <= 24'd00633967;
                12'd1519: logsin <= 24'd00634706;
                12'd1520: logsin <= 24'd00635445;
                12'd1521: logsin <= 24'd00636185;
                12'd1522: logsin <= 24'd00636924;
                12'd1523: logsin <= 24'd00637664;
                12'd1524: logsin <= 24'd00638404;
                12'd1525: logsin <= 24'd00639144;
                12'd1526: logsin <= 24'd00639885;
                12'd1527: logsin <= 24'd00640626;
                12'd1528: logsin <= 24'd00641367;
                12'd1529: logsin <= 24'd00642108;
                12'd1530: logsin <= 24'd00642849;
                12'd1531: logsin <= 24'd00643591;
                12'd1532: logsin <= 24'd00644333;
                12'd1533: logsin <= 24'd00645075;
                12'd1534: logsin <= 24'd00645818;
                12'd1535: logsin <= 24'd00646560;
                12'd1536: logsin <= 24'd00647303;
                12'd1537: logsin <= 24'd00648046;
                12'd1538: logsin <= 24'd00648790;
                12'd1539: logsin <= 24'd00649533;
                12'd1540: logsin <= 24'd00650277;
                12'd1541: logsin <= 24'd00651021;
                12'd1542: logsin <= 24'd00651766;
                12'd1543: logsin <= 24'd00652510;
                12'd1544: logsin <= 24'd00653255;
                12'd1545: logsin <= 24'd00654000;
                12'd1546: logsin <= 24'd00654745;
                12'd1547: logsin <= 24'd00655491;
                12'd1548: logsin <= 24'd00656237;
                12'd1549: logsin <= 24'd00656982;
                12'd1550: logsin <= 24'd00657729;
                12'd1551: logsin <= 24'd00658475;
                12'd1552: logsin <= 24'd00659222;
                12'd1553: logsin <= 24'd00659969;
                12'd1554: logsin <= 24'd00660716;
                12'd1555: logsin <= 24'd00661463;
                12'd1556: logsin <= 24'd00662211;
                12'd1557: logsin <= 24'd00662958;
                12'd1558: logsin <= 24'd00663706;
                12'd1559: logsin <= 24'd00664455;
                12'd1560: logsin <= 24'd00665203;
                12'd1561: logsin <= 24'd00665952;
                12'd1562: logsin <= 24'd00666701;
                12'd1563: logsin <= 24'd00667450;
                12'd1564: logsin <= 24'd00668199;
                12'd1565: logsin <= 24'd00668949;
                12'd1566: logsin <= 24'd00669698;
                12'd1567: logsin <= 24'd00670448;
                12'd1568: logsin <= 24'd00671199;
                12'd1569: logsin <= 24'd00671949;
                12'd1570: logsin <= 24'd00672700;
                12'd1571: logsin <= 24'd00673451;
                12'd1572: logsin <= 24'd00674202;
                12'd1573: logsin <= 24'd00674953;
                12'd1574: logsin <= 24'd00675705;
                12'd1575: logsin <= 24'd00676457;
                12'd1576: logsin <= 24'd00677209;
                12'd1577: logsin <= 24'd00677961;
                12'd1578: logsin <= 24'd00678713;
                12'd1579: logsin <= 24'd00679466;
                12'd1580: logsin <= 24'd00680219;
                12'd1581: logsin <= 24'd00680972;
                12'd1582: logsin <= 24'd00681725;
                12'd1583: logsin <= 24'd00682479;
                12'd1584: logsin <= 24'd00683233;
                12'd1585: logsin <= 24'd00683986;
                12'd1586: logsin <= 24'd00684741;
                12'd1587: logsin <= 24'd00685495;
                12'd1588: logsin <= 24'd00686250;
                12'd1589: logsin <= 24'd00687004;
                12'd1590: logsin <= 24'd00687760;
                12'd1591: logsin <= 24'd00688515;
                12'd1592: logsin <= 24'd00689270;
                12'd1593: logsin <= 24'd00690026;
                12'd1594: logsin <= 24'd00690782;
                12'd1595: logsin <= 24'd00691538;
                12'd1596: logsin <= 24'd00692294;
                12'd1597: logsin <= 24'd00693051;
                12'd1598: logsin <= 24'd00693807;
                12'd1599: logsin <= 24'd00694564;
                12'd1600: logsin <= 24'd00695321;
                12'd1601: logsin <= 24'd00696079;
                12'd1602: logsin <= 24'd00696836;
                12'd1603: logsin <= 24'd00697594;
                12'd1604: logsin <= 24'd00698352;
                12'd1605: logsin <= 24'd00699110;
                12'd1606: logsin <= 24'd00699869;
                12'd1607: logsin <= 24'd00700627;
                12'd1608: logsin <= 24'd00701386;
                12'd1609: logsin <= 24'd00702145;
                12'd1610: logsin <= 24'd00702904;
                12'd1611: logsin <= 24'd00703663;
                12'd1612: logsin <= 24'd00704423;
                12'd1613: logsin <= 24'd00705183;
                12'd1614: logsin <= 24'd00705943;
                12'd1615: logsin <= 24'd00706703;
                12'd1616: logsin <= 24'd00707463;
                12'd1617: logsin <= 24'd00708224;
                12'd1618: logsin <= 24'd00708985;
                12'd1619: logsin <= 24'd00709746;
                12'd1620: logsin <= 24'd00710507;
                12'd1621: logsin <= 24'd00711268;
                12'd1622: logsin <= 24'd00712030;
                12'd1623: logsin <= 24'd00712792;
                12'd1624: logsin <= 24'd00713554;
                12'd1625: logsin <= 24'd00714316;
                12'd1626: logsin <= 24'd00715078;
                12'd1627: logsin <= 24'd00715841;
                12'd1628: logsin <= 24'd00716604;
                12'd1629: logsin <= 24'd00717367;
                12'd1630: logsin <= 24'd00718130;
                12'd1631: logsin <= 24'd00718893;
                12'd1632: logsin <= 24'd00719657;
                12'd1633: logsin <= 24'd00720421;
                12'd1634: logsin <= 24'd00721185;
                12'd1635: logsin <= 24'd00721949;
                12'd1636: logsin <= 24'd00722713;
                12'd1637: logsin <= 24'd00723478;
                12'd1638: logsin <= 24'd00724242;
                12'd1639: logsin <= 24'd00725007;
                12'd1640: logsin <= 24'd00725772;
                12'd1641: logsin <= 24'd00726538;
                12'd1642: logsin <= 24'd00727303;
                12'd1643: logsin <= 24'd00728069;
                12'd1644: logsin <= 24'd00728835;
                12'd1645: logsin <= 24'd00729601;
                12'd1646: logsin <= 24'd00730367;
                12'd1647: logsin <= 24'd00731133;
                12'd1648: logsin <= 24'd00731900;
                12'd1649: logsin <= 24'd00732667;
                12'd1650: logsin <= 24'd00733434;
                12'd1651: logsin <= 24'd00734201;
                12'd1652: logsin <= 24'd00734968;
                12'd1653: logsin <= 24'd00735736;
                12'd1654: logsin <= 24'd00736503;
                12'd1655: logsin <= 24'd00737271;
                12'd1656: logsin <= 24'd00738039;
                12'd1657: logsin <= 24'd00738808;
                12'd1658: logsin <= 24'd00739576;
                12'd1659: logsin <= 24'd00740345;
                12'd1660: logsin <= 24'd00741113;
                12'd1661: logsin <= 24'd00741882;
                12'd1662: logsin <= 24'd00742652;
                12'd1663: logsin <= 24'd00743421;
                12'd1664: logsin <= 24'd00744190;
                12'd1665: logsin <= 24'd00744960;
                12'd1666: logsin <= 24'd00745730;
                12'd1667: logsin <= 24'd00746500;
                12'd1668: logsin <= 24'd00747270;
                12'd1669: logsin <= 24'd00748041;
                12'd1670: logsin <= 24'd00748811;
                12'd1671: logsin <= 24'd00749582;
                12'd1672: logsin <= 24'd00750353;
                12'd1673: logsin <= 24'd00751124;
                12'd1674: logsin <= 24'd00751896;
                12'd1675: logsin <= 24'd00752667;
                12'd1676: logsin <= 24'd00753439;
                12'd1677: logsin <= 24'd00754210;
                12'd1678: logsin <= 24'd00754982;
                12'd1679: logsin <= 24'd00755755;
                12'd1680: logsin <= 24'd00756527;
                12'd1681: logsin <= 24'd00757299;
                12'd1682: logsin <= 24'd00758072;
                12'd1683: logsin <= 24'd00758845;
                12'd1684: logsin <= 24'd00759618;
                12'd1685: logsin <= 24'd00760391;
                12'd1686: logsin <= 24'd00761165;
                12'd1687: logsin <= 24'd00761938;
                12'd1688: logsin <= 24'd00762712;
                12'd1689: logsin <= 24'd00763486;
                12'd1690: logsin <= 24'd00764260;
                12'd1691: logsin <= 24'd00765034;
                12'd1692: logsin <= 24'd00765808;
                12'd1693: logsin <= 24'd00766583;
                12'd1694: logsin <= 24'd00767358;
                12'd1695: logsin <= 24'd00768132;
                12'd1696: logsin <= 24'd00768907;
                12'd1697: logsin <= 24'd00769683;
                12'd1698: logsin <= 24'd00770458;
                12'd1699: logsin <= 24'd00771233;
                12'd1700: logsin <= 24'd00772009;
                12'd1701: logsin <= 24'd00772785;
                12'd1702: logsin <= 24'd00773561;
                12'd1703: logsin <= 24'd00774337;
                12'd1704: logsin <= 24'd00775114;
                12'd1705: logsin <= 24'd00775890;
                12'd1706: logsin <= 24'd00776667;
                12'd1707: logsin <= 24'd00777444;
                12'd1708: logsin <= 24'd00778220;
                12'd1709: logsin <= 24'd00778998;
                12'd1710: logsin <= 24'd00779775;
                12'd1711: logsin <= 24'd00780552;
                12'd1712: logsin <= 24'd00781330;
                12'd1713: logsin <= 24'd00782108;
                12'd1714: logsin <= 24'd00782886;
                12'd1715: logsin <= 24'd00783664;
                12'd1716: logsin <= 24'd00784442;
                12'd1717: logsin <= 24'd00785220;
                12'd1718: logsin <= 24'd00785999;
                12'd1719: logsin <= 24'd00786778;
                12'd1720: logsin <= 24'd00787556;
                12'd1721: logsin <= 24'd00788335;
                12'd1722: logsin <= 24'd00789115;
                12'd1723: logsin <= 24'd00789894;
                12'd1724: logsin <= 24'd00790673;
                12'd1725: logsin <= 24'd00791453;
                12'd1726: logsin <= 24'd00792233;
                12'd1727: logsin <= 24'd00793013;
                12'd1728: logsin <= 24'd00793793;
                12'd1729: logsin <= 24'd00794573;
                12'd1730: logsin <= 24'd00795353;
                12'd1731: logsin <= 24'd00796134;
                12'd1732: logsin <= 24'd00796915;
                12'd1733: logsin <= 24'd00797695;
                12'd1734: logsin <= 24'd00798476;
                12'd1735: logsin <= 24'd00799257;
                12'd1736: logsin <= 24'd00800039;
                12'd1737: logsin <= 24'd00800820;
                12'd1738: logsin <= 24'd00801602;
                12'd1739: logsin <= 24'd00802383;
                12'd1740: logsin <= 24'd00803165;
                12'd1741: logsin <= 24'd00803947;
                12'd1742: logsin <= 24'd00804729;
                12'd1743: logsin <= 24'd00805512;
                12'd1744: logsin <= 24'd00806294;
                12'd1745: logsin <= 24'd00807077;
                12'd1746: logsin <= 24'd00807859;
                12'd1747: logsin <= 24'd00808642;
                12'd1748: logsin <= 24'd00809425;
                12'd1749: logsin <= 24'd00810208;
                12'd1750: logsin <= 24'd00810991;
                12'd1751: logsin <= 24'd00811775;
                12'd1752: logsin <= 24'd00812558;
                12'd1753: logsin <= 24'd00813342;
                12'd1754: logsin <= 24'd00814126;
                12'd1755: logsin <= 24'd00814910;
                12'd1756: logsin <= 24'd00815694;
                12'd1757: logsin <= 24'd00816478;
                12'd1758: logsin <= 24'd00817263;
                12'd1759: logsin <= 24'd00818047;
                12'd1760: logsin <= 24'd00818832;
                12'd1761: logsin <= 24'd00819616;
                12'd1762: logsin <= 24'd00820401;
                12'd1763: logsin <= 24'd00821186;
                12'd1764: logsin <= 24'd00821972;
                12'd1765: logsin <= 24'd00822757;
                12'd1766: logsin <= 24'd00823542;
                12'd1767: logsin <= 24'd00824328;
                12'd1768: logsin <= 24'd00825114;
                12'd1769: logsin <= 24'd00825899;
                12'd1770: logsin <= 24'd00826685;
                12'd1771: logsin <= 24'd00827472;
                12'd1772: logsin <= 24'd00828258;
                12'd1773: logsin <= 24'd00829044;
                12'd1774: logsin <= 24'd00829831;
                12'd1775: logsin <= 24'd00830617;
                12'd1776: logsin <= 24'd00831404;
                12'd1777: logsin <= 24'd00832191;
                12'd1778: logsin <= 24'd00832978;
                12'd1779: logsin <= 24'd00833765;
                12'd1780: logsin <= 24'd00834552;
                12'd1781: logsin <= 24'd00835340;
                12'd1782: logsin <= 24'd00836127;
                12'd1783: logsin <= 24'd00836915;
                12'd1784: logsin <= 24'd00837703;
                12'd1785: logsin <= 24'd00838490;
                12'd1786: logsin <= 24'd00839278;
                12'd1787: logsin <= 24'd00840067;
                12'd1788: logsin <= 24'd00840855;
                12'd1789: logsin <= 24'd00841643;
                12'd1790: logsin <= 24'd00842432;
                12'd1791: logsin <= 24'd00843220;
                12'd1792: logsin <= 24'd00844009;
                12'd1793: logsin <= 24'd00844798;
                12'd1794: logsin <= 24'd00845587;
                12'd1795: logsin <= 24'd00846376;
                12'd1796: logsin <= 24'd00847165;
                12'd1797: logsin <= 24'd00847954;
                12'd1798: logsin <= 24'd00848744;
                12'd1799: logsin <= 24'd00849533;
                12'd1800: logsin <= 24'd00850323;
                12'd1801: logsin <= 24'd00851113;
                12'd1802: logsin <= 24'd00851903;
                12'd1803: logsin <= 24'd00852693;
                12'd1804: logsin <= 24'd00853483;
                12'd1805: logsin <= 24'd00854273;
                12'd1806: logsin <= 24'd00855064;
                12'd1807: logsin <= 24'd00855854;
                12'd1808: logsin <= 24'd00856645;
                12'd1809: logsin <= 24'd00857435;
                12'd1810: logsin <= 24'd00858226;
                12'd1811: logsin <= 24'd00859017;
                12'd1812: logsin <= 24'd00859808;
                12'd1813: logsin <= 24'd00860599;
                12'd1814: logsin <= 24'd00861391;
                12'd1815: logsin <= 24'd00862182;
                12'd1816: logsin <= 24'd00862974;
                12'd1817: logsin <= 24'd00863765;
                12'd1818: logsin <= 24'd00864557;
                12'd1819: logsin <= 24'd00865349;
                12'd1820: logsin <= 24'd00866141;
                12'd1821: logsin <= 24'd00866933;
                12'd1822: logsin <= 24'd00867725;
                12'd1823: logsin <= 24'd00868517;
                12'd1824: logsin <= 24'd00869309;
                12'd1825: logsin <= 24'd00870102;
                12'd1826: logsin <= 24'd00870894;
                12'd1827: logsin <= 24'd00871687;
                12'd1828: logsin <= 24'd00872480;
                12'd1829: logsin <= 24'd00873273;
                12'd1830: logsin <= 24'd00874066;
                12'd1831: logsin <= 24'd00874859;
                12'd1832: logsin <= 24'd00875652;
                12'd1833: logsin <= 24'd00876445;
                12'd1834: logsin <= 24'd00877239;
                12'd1835: logsin <= 24'd00878032;
                12'd1836: logsin <= 24'd00878826;
                12'd1837: logsin <= 24'd00879620;
                12'd1838: logsin <= 24'd00880413;
                12'd1839: logsin <= 24'd00881207;
                12'd1840: logsin <= 24'd00882001;
                12'd1841: logsin <= 24'd00882795;
                12'd1842: logsin <= 24'd00883589;
                12'd1843: logsin <= 24'd00884384;
                12'd1844: logsin <= 24'd00885178;
                12'd1845: logsin <= 24'd00885973;
                12'd1846: logsin <= 24'd00886767;
                12'd1847: logsin <= 24'd00887562;
                12'd1848: logsin <= 24'd00888357;
                12'd1849: logsin <= 24'd00889151;
                12'd1850: logsin <= 24'd00889946;
                12'd1851: logsin <= 24'd00890741;
                12'd1852: logsin <= 24'd00891537;
                12'd1853: logsin <= 24'd00892332;
                12'd1854: logsin <= 24'd00893127;
                12'd1855: logsin <= 24'd00893922;
                12'd1856: logsin <= 24'd00894718;
                12'd1857: logsin <= 24'd00895514;
                12'd1858: logsin <= 24'd00896309;
                12'd1859: logsin <= 24'd00897105;
                12'd1860: logsin <= 24'd00897901;
                12'd1861: logsin <= 24'd00898697;
                12'd1862: logsin <= 24'd00899493;
                12'd1863: logsin <= 24'd00900289;
                12'd1864: logsin <= 24'd00901085;
                12'd1865: logsin <= 24'd00901881;
                12'd1866: logsin <= 24'd00902678;
                12'd1867: logsin <= 24'd00903474;
                12'd1868: logsin <= 24'd00904271;
                12'd1869: logsin <= 24'd00905067;
                12'd1870: logsin <= 24'd00905864;
                12'd1871: logsin <= 24'd00906661;
                12'd1872: logsin <= 24'd00907458;
                12'd1873: logsin <= 24'd00908255;
                12'd1874: logsin <= 24'd00909052;
                12'd1875: logsin <= 24'd00909849;
                12'd1876: logsin <= 24'd00910646;
                12'd1877: logsin <= 24'd00911444;
                12'd1878: logsin <= 24'd00912241;
                12'd1879: logsin <= 24'd00913038;
                12'd1880: logsin <= 24'd00913836;
                12'd1881: logsin <= 24'd00914634;
                12'd1882: logsin <= 24'd00915431;
                12'd1883: logsin <= 24'd00916229;
                12'd1884: logsin <= 24'd00917027;
                12'd1885: logsin <= 24'd00917825;
                12'd1886: logsin <= 24'd00918623;
                12'd1887: logsin <= 24'd00919421;
                12'd1888: logsin <= 24'd00920219;
                12'd1889: logsin <= 24'd00921017;
                12'd1890: logsin <= 24'd00921816;
                12'd1891: logsin <= 24'd00922614;
                12'd1892: logsin <= 24'd00923413;
                12'd1893: logsin <= 24'd00924211;
                12'd1894: logsin <= 24'd00925010;
                12'd1895: logsin <= 24'd00925808;
                12'd1896: logsin <= 24'd00926607;
                12'd1897: logsin <= 24'd00927406;
                12'd1898: logsin <= 24'd00928205;
                12'd1899: logsin <= 24'd00929004;
                12'd1900: logsin <= 24'd00929803;
                12'd1901: logsin <= 24'd00930602;
                12'd1902: logsin <= 24'd00931401;
                12'd1903: logsin <= 24'd00932200;
                12'd1904: logsin <= 24'd00933000;
                12'd1905: logsin <= 24'd00933799;
                12'd1906: logsin <= 24'd00934598;
                12'd1907: logsin <= 24'd00935398;
                12'd1908: logsin <= 24'd00936198;
                12'd1909: logsin <= 24'd00936997;
                12'd1910: logsin <= 24'd00937797;
                12'd1911: logsin <= 24'd00938597;
                12'd1912: logsin <= 24'd00939397;
                12'd1913: logsin <= 24'd00940196;
                12'd1914: logsin <= 24'd00940996;
                12'd1915: logsin <= 24'd00941796;
                12'd1916: logsin <= 24'd00942597;
                12'd1917: logsin <= 24'd00943397;
                12'd1918: logsin <= 24'd00944197;
                12'd1919: logsin <= 24'd00944997;
                12'd1920: logsin <= 24'd00945798;
                12'd1921: logsin <= 24'd00946598;
                12'd1922: logsin <= 24'd00947398;
                12'd1923: logsin <= 24'd00948199;
                12'd1924: logsin <= 24'd00949000;
                12'd1925: logsin <= 24'd00949800;
                12'd1926: logsin <= 24'd00950601;
                12'd1927: logsin <= 24'd00951402;
                12'd1928: logsin <= 24'd00952202;
                12'd1929: logsin <= 24'd00953003;
                12'd1930: logsin <= 24'd00953804;
                12'd1931: logsin <= 24'd00954605;
                12'd1932: logsin <= 24'd00955406;
                12'd1933: logsin <= 24'd00956207;
                12'd1934: logsin <= 24'd00957009;
                12'd1935: logsin <= 24'd00957810;
                12'd1936: logsin <= 24'd00958611;
                12'd1937: logsin <= 24'd00959412;
                12'd1938: logsin <= 24'd00960214;
                12'd1939: logsin <= 24'd00961015;
                12'd1940: logsin <= 24'd00961817;
                12'd1941: logsin <= 24'd00962618;
                12'd1942: logsin <= 24'd00963420;
                12'd1943: logsin <= 24'd00964221;
                12'd1944: logsin <= 24'd00965023;
                12'd1945: logsin <= 24'd00965825;
                12'd1946: logsin <= 24'd00966626;
                12'd1947: logsin <= 24'd00967428;
                12'd1948: logsin <= 24'd00968230;
                12'd1949: logsin <= 24'd00969032;
                12'd1950: logsin <= 24'd00969834;
                12'd1951: logsin <= 24'd00970636;
                12'd1952: logsin <= 24'd00971438;
                12'd1953: logsin <= 24'd00972240;
                12'd1954: logsin <= 24'd00973042;
                12'd1955: logsin <= 24'd00973844;
                12'd1956: logsin <= 24'd00974647;
                12'd1957: logsin <= 24'd00975449;
                12'd1958: logsin <= 24'd00976251;
                12'd1959: logsin <= 24'd00977054;
                12'd1960: logsin <= 24'd00977856;
                12'd1961: logsin <= 24'd00978658;
                12'd1962: logsin <= 24'd00979461;
                12'd1963: logsin <= 24'd00980263;
                12'd1964: logsin <= 24'd00981066;
                12'd1965: logsin <= 24'd00981869;
                12'd1966: logsin <= 24'd00982671;
                12'd1967: logsin <= 24'd00983474;
                12'd1968: logsin <= 24'd00984277;
                12'd1969: logsin <= 24'd00985079;
                12'd1970: logsin <= 24'd00985882;
                12'd1971: logsin <= 24'd00986685;
                12'd1972: logsin <= 24'd00987488;
                12'd1973: logsin <= 24'd00988291;
                12'd1974: logsin <= 24'd00989094;
                12'd1975: logsin <= 24'd00989897;
                12'd1976: logsin <= 24'd00990700;
                12'd1977: logsin <= 24'd00991503;
                12'd1978: logsin <= 24'd00992306;
                12'd1979: logsin <= 24'd00993109;
                12'd1980: logsin <= 24'd00993912;
                12'd1981: logsin <= 24'd00994715;
                12'd1982: logsin <= 24'd00995518;
                12'd1983: logsin <= 24'd00996322;
                12'd1984: logsin <= 24'd00997125;
                12'd1985: logsin <= 24'd00997928;
                12'd1986: logsin <= 24'd00998731;
                12'd1987: logsin <= 24'd00999535;
                12'd1988: logsin <= 24'd01000338;
                12'd1989: logsin <= 24'd01001142;
                12'd1990: logsin <= 24'd01001945;
                12'd1991: logsin <= 24'd01002748;
                12'd1992: logsin <= 24'd01003552;
                12'd1993: logsin <= 24'd01004355;
                12'd1994: logsin <= 24'd01005159;
                12'd1995: logsin <= 24'd01005963;
                12'd1996: logsin <= 24'd01006766;
                12'd1997: logsin <= 24'd01007570;
                12'd1998: logsin <= 24'd01008373;
                12'd1999: logsin <= 24'd01009177;
                12'd2000: logsin <= 24'd01009981;
                12'd2001: logsin <= 24'd01010785;
                12'd2002: logsin <= 24'd01011588;
                12'd2003: logsin <= 24'd01012392;
                12'd2004: logsin <= 24'd01013196;
                12'd2005: logsin <= 24'd01014000;
                12'd2006: logsin <= 24'd01014803;
                12'd2007: logsin <= 24'd01015607;
                12'd2008: logsin <= 24'd01016411;
                12'd2009: logsin <= 24'd01017215;
                12'd2010: logsin <= 24'd01018019;
                12'd2011: logsin <= 24'd01018823;
                12'd2012: logsin <= 24'd01019627;
                12'd2013: logsin <= 24'd01020431;
                12'd2014: logsin <= 24'd01021235;
                12'd2015: logsin <= 24'd01022039;
                12'd2016: logsin <= 24'd01022843;
                12'd2017: logsin <= 24'd01023647;
                12'd2018: logsin <= 24'd01024451;
                12'd2019: logsin <= 24'd01025255;
                12'd2020: logsin <= 24'd01026059;
                12'd2021: logsin <= 24'd01026863;
                12'd2022: logsin <= 24'd01027667;
                12'd2023: logsin <= 24'd01028471;
                12'd2024: logsin <= 24'd01029275;
                12'd2025: logsin <= 24'd01030079;
                12'd2026: logsin <= 24'd01030883;
                12'd2027: logsin <= 24'd01031688;
                12'd2028: logsin <= 24'd01032492;
                12'd2029: logsin <= 24'd01033296;
                12'd2030: logsin <= 24'd01034100;
                12'd2031: logsin <= 24'd01034904;
                12'd2032: logsin <= 24'd01035708;
                12'd2033: logsin <= 24'd01036513;
                12'd2034: logsin <= 24'd01037317;
                12'd2035: logsin <= 24'd01038121;
                12'd2036: logsin <= 24'd01038925;
                12'd2037: logsin <= 24'd01039729;
                12'd2038: logsin <= 24'd01040534;
                12'd2039: logsin <= 24'd01041338;
                12'd2040: logsin <= 24'd01042142;
                12'd2041: logsin <= 24'd01042946;
                12'd2042: logsin <= 24'd01043751;
                12'd2043: logsin <= 24'd01044555;
                12'd2044: logsin <= 24'd01045359;
                12'd2045: logsin <= 24'd01046163;
                12'd2046: logsin <= 24'd01046968;
                12'd2047: logsin <= 24'd01047772;
                12'd2048: logsin <= 24'd01048576;
                12'd2049: logsin <= 24'd01049380;
                12'd2050: logsin <= 24'd01050184;
                12'd2051: logsin <= 24'd01050989;
                12'd2052: logsin <= 24'd01051793;
                12'd2053: logsin <= 24'd01052597;
                12'd2054: logsin <= 24'd01053401;
                12'd2055: logsin <= 24'd01054206;
                12'd2056: logsin <= 24'd01055010;
                12'd2057: logsin <= 24'd01055814;
                12'd2058: logsin <= 24'd01056618;
                12'd2059: logsin <= 24'd01057423;
                12'd2060: logsin <= 24'd01058227;
                12'd2061: logsin <= 24'd01059031;
                12'd2062: logsin <= 24'd01059835;
                12'd2063: logsin <= 24'd01060639;
                12'd2064: logsin <= 24'd01061444;
                12'd2065: logsin <= 24'd01062248;
                12'd2066: logsin <= 24'd01063052;
                12'd2067: logsin <= 24'd01063856;
                12'd2068: logsin <= 24'd01064660;
                12'd2069: logsin <= 24'd01065464;
                12'd2070: logsin <= 24'd01066269;
                12'd2071: logsin <= 24'd01067073;
                12'd2072: logsin <= 24'd01067877;
                12'd2073: logsin <= 24'd01068681;
                12'd2074: logsin <= 24'd01069485;
                12'd2075: logsin <= 24'd01070289;
                12'd2076: logsin <= 24'd01071093;
                12'd2077: logsin <= 24'd01071897;
                12'd2078: logsin <= 24'd01072701;
                12'd2079: logsin <= 24'd01073505;
                12'd2080: logsin <= 24'd01074309;
                12'd2081: logsin <= 24'd01075113;
                12'd2082: logsin <= 24'd01075917;
                12'd2083: logsin <= 24'd01076721;
                12'd2084: logsin <= 24'd01077525;
                12'd2085: logsin <= 24'd01078329;
                12'd2086: logsin <= 24'd01079133;
                12'd2087: logsin <= 24'd01079937;
                12'd2088: logsin <= 24'd01080741;
                12'd2089: logsin <= 24'd01081545;
                12'd2090: logsin <= 24'd01082349;
                12'd2091: logsin <= 24'd01083152;
                12'd2092: logsin <= 24'd01083956;
                12'd2093: logsin <= 24'd01084760;
                12'd2094: logsin <= 24'd01085564;
                12'd2095: logsin <= 24'd01086367;
                12'd2096: logsin <= 24'd01087171;
                12'd2097: logsin <= 24'd01087975;
                12'd2098: logsin <= 24'd01088779;
                12'd2099: logsin <= 24'd01089582;
                12'd2100: logsin <= 24'd01090386;
                12'd2101: logsin <= 24'd01091189;
                12'd2102: logsin <= 24'd01091993;
                12'd2103: logsin <= 24'd01092797;
                12'd2104: logsin <= 24'd01093600;
                12'd2105: logsin <= 24'd01094404;
                12'd2106: logsin <= 24'd01095207;
                12'd2107: logsin <= 24'd01096010;
                12'd2108: logsin <= 24'd01096814;
                12'd2109: logsin <= 24'd01097617;
                12'd2110: logsin <= 24'd01098421;
                12'd2111: logsin <= 24'd01099224;
                12'd2112: logsin <= 24'd01100027;
                12'd2113: logsin <= 24'd01100830;
                12'd2114: logsin <= 24'd01101634;
                12'd2115: logsin <= 24'd01102437;
                12'd2116: logsin <= 24'd01103240;
                12'd2117: logsin <= 24'd01104043;
                12'd2118: logsin <= 24'd01104846;
                12'd2119: logsin <= 24'd01105649;
                12'd2120: logsin <= 24'd01106452;
                12'd2121: logsin <= 24'd01107255;
                12'd2122: logsin <= 24'd01108058;
                12'd2123: logsin <= 24'd01108861;
                12'd2124: logsin <= 24'd01109664;
                12'd2125: logsin <= 24'd01110467;
                12'd2126: logsin <= 24'd01111270;
                12'd2127: logsin <= 24'd01112073;
                12'd2128: logsin <= 24'd01112875;
                12'd2129: logsin <= 24'd01113678;
                12'd2130: logsin <= 24'd01114481;
                12'd2131: logsin <= 24'd01115283;
                12'd2132: logsin <= 24'd01116086;
                12'd2133: logsin <= 24'd01116889;
                12'd2134: logsin <= 24'd01117691;
                12'd2135: logsin <= 24'd01118494;
                12'd2136: logsin <= 24'd01119296;
                12'd2137: logsin <= 24'd01120098;
                12'd2138: logsin <= 24'd01120901;
                12'd2139: logsin <= 24'd01121703;
                12'd2140: logsin <= 24'd01122505;
                12'd2141: logsin <= 24'd01123308;
                12'd2142: logsin <= 24'd01124110;
                12'd2143: logsin <= 24'd01124912;
                12'd2144: logsin <= 24'd01125714;
                12'd2145: logsin <= 24'd01126516;
                12'd2146: logsin <= 24'd01127318;
                12'd2147: logsin <= 24'd01128120;
                12'd2148: logsin <= 24'd01128922;
                12'd2149: logsin <= 24'd01129724;
                12'd2150: logsin <= 24'd01130526;
                12'd2151: logsin <= 24'd01131327;
                12'd2152: logsin <= 24'd01132129;
                12'd2153: logsin <= 24'd01132931;
                12'd2154: logsin <= 24'd01133732;
                12'd2155: logsin <= 24'd01134534;
                12'd2156: logsin <= 24'd01135335;
                12'd2157: logsin <= 24'd01136137;
                12'd2158: logsin <= 24'd01136938;
                12'd2159: logsin <= 24'd01137740;
                12'd2160: logsin <= 24'd01138541;
                12'd2161: logsin <= 24'd01139342;
                12'd2162: logsin <= 24'd01140143;
                12'd2163: logsin <= 24'd01140945;
                12'd2164: logsin <= 24'd01141746;
                12'd2165: logsin <= 24'd01142547;
                12'd2166: logsin <= 24'd01143348;
                12'd2167: logsin <= 24'd01144149;
                12'd2168: logsin <= 24'd01144950;
                12'd2169: logsin <= 24'd01145750;
                12'd2170: logsin <= 24'd01146551;
                12'd2171: logsin <= 24'd01147352;
                12'd2172: logsin <= 24'd01148152;
                12'd2173: logsin <= 24'd01148953;
                12'd2174: logsin <= 24'd01149754;
                12'd2175: logsin <= 24'd01150554;
                12'd2176: logsin <= 24'd01151354;
                12'd2177: logsin <= 24'd01152155;
                12'd2178: logsin <= 24'd01152955;
                12'd2179: logsin <= 24'd01153755;
                12'd2180: logsin <= 24'd01154555;
                12'd2181: logsin <= 24'd01155356;
                12'd2182: logsin <= 24'd01156156;
                12'd2183: logsin <= 24'd01156956;
                12'd2184: logsin <= 24'd01157755;
                12'd2185: logsin <= 24'd01158555;
                12'd2186: logsin <= 24'd01159355;
                12'd2187: logsin <= 24'd01160155;
                12'd2188: logsin <= 24'd01160954;
                12'd2189: logsin <= 24'd01161754;
                12'd2190: logsin <= 24'd01162554;
                12'd2191: logsin <= 24'd01163353;
                12'd2192: logsin <= 24'd01164152;
                12'd2193: logsin <= 24'd01164952;
                12'd2194: logsin <= 24'd01165751;
                12'd2195: logsin <= 24'd01166550;
                12'd2196: logsin <= 24'd01167349;
                12'd2197: logsin <= 24'd01168148;
                12'd2198: logsin <= 24'd01168947;
                12'd2199: logsin <= 24'd01169746;
                12'd2200: logsin <= 24'd01170545;
                12'd2201: logsin <= 24'd01171344;
                12'd2202: logsin <= 24'd01172142;
                12'd2203: logsin <= 24'd01172941;
                12'd2204: logsin <= 24'd01173739;
                12'd2205: logsin <= 24'd01174538;
                12'd2206: logsin <= 24'd01175336;
                12'd2207: logsin <= 24'd01176135;
                12'd2208: logsin <= 24'd01176933;
                12'd2209: logsin <= 24'd01177731;
                12'd2210: logsin <= 24'd01178529;
                12'd2211: logsin <= 24'd01179327;
                12'd2212: logsin <= 24'd01180125;
                12'd2213: logsin <= 24'd01180923;
                12'd2214: logsin <= 24'd01181721;
                12'd2215: logsin <= 24'd01182518;
                12'd2216: logsin <= 24'd01183316;
                12'd2217: logsin <= 24'd01184114;
                12'd2218: logsin <= 24'd01184911;
                12'd2219: logsin <= 24'd01185708;
                12'd2220: logsin <= 24'd01186506;
                12'd2221: logsin <= 24'd01187303;
                12'd2222: logsin <= 24'd01188100;
                12'd2223: logsin <= 24'd01188897;
                12'd2224: logsin <= 24'd01189694;
                12'd2225: logsin <= 24'd01190491;
                12'd2226: logsin <= 24'd01191288;
                12'd2227: logsin <= 24'd01192085;
                12'd2228: logsin <= 24'd01192881;
                12'd2229: logsin <= 24'd01193678;
                12'd2230: logsin <= 24'd01194474;
                12'd2231: logsin <= 24'd01195271;
                12'd2232: logsin <= 24'd01196067;
                12'd2233: logsin <= 24'd01196863;
                12'd2234: logsin <= 24'd01197659;
                12'd2235: logsin <= 24'd01198455;
                12'd2236: logsin <= 24'd01199251;
                12'd2237: logsin <= 24'd01200047;
                12'd2238: logsin <= 24'd01200843;
                12'd2239: logsin <= 24'd01201638;
                12'd2240: logsin <= 24'd01202434;
                12'd2241: logsin <= 24'd01203230;
                12'd2242: logsin <= 24'd01204025;
                12'd2243: logsin <= 24'd01204820;
                12'd2244: logsin <= 24'd01205615;
                12'd2245: logsin <= 24'd01206411;
                12'd2246: logsin <= 24'd01207206;
                12'd2247: logsin <= 24'd01208001;
                12'd2248: logsin <= 24'd01208795;
                12'd2249: logsin <= 24'd01209590;
                12'd2250: logsin <= 24'd01210385;
                12'd2251: logsin <= 24'd01211179;
                12'd2252: logsin <= 24'd01211974;
                12'd2253: logsin <= 24'd01212768;
                12'd2254: logsin <= 24'd01213563;
                12'd2255: logsin <= 24'd01214357;
                12'd2256: logsin <= 24'd01215151;
                12'd2257: logsin <= 24'd01215945;
                12'd2258: logsin <= 24'd01216739;
                12'd2259: logsin <= 24'd01217532;
                12'd2260: logsin <= 24'd01218326;
                12'd2261: logsin <= 24'd01219120;
                12'd2262: logsin <= 24'd01219913;
                12'd2263: logsin <= 24'd01220707;
                12'd2264: logsin <= 24'd01221500;
                12'd2265: logsin <= 24'd01222293;
                12'd2266: logsin <= 24'd01223086;
                12'd2267: logsin <= 24'd01223879;
                12'd2268: logsin <= 24'd01224672;
                12'd2269: logsin <= 24'd01225465;
                12'd2270: logsin <= 24'd01226258;
                12'd2271: logsin <= 24'd01227050;
                12'd2272: logsin <= 24'd01227843;
                12'd2273: logsin <= 24'd01228635;
                12'd2274: logsin <= 24'd01229427;
                12'd2275: logsin <= 24'd01230219;
                12'd2276: logsin <= 24'd01231011;
                12'd2277: logsin <= 24'd01231803;
                12'd2278: logsin <= 24'd01232595;
                12'd2279: logsin <= 24'd01233387;
                12'd2280: logsin <= 24'd01234178;
                12'd2281: logsin <= 24'd01234970;
                12'd2282: logsin <= 24'd01235761;
                12'd2283: logsin <= 24'd01236553;
                12'd2284: logsin <= 24'd01237344;
                12'd2285: logsin <= 24'd01238135;
                12'd2286: logsin <= 24'd01238926;
                12'd2287: logsin <= 24'd01239717;
                12'd2288: logsin <= 24'd01240507;
                12'd2289: logsin <= 24'd01241298;
                12'd2290: logsin <= 24'd01242088;
                12'd2291: logsin <= 24'd01242879;
                12'd2292: logsin <= 24'd01243669;
                12'd2293: logsin <= 24'd01244459;
                12'd2294: logsin <= 24'd01245249;
                12'd2295: logsin <= 24'd01246039;
                12'd2296: logsin <= 24'd01246829;
                12'd2297: logsin <= 24'd01247619;
                12'd2298: logsin <= 24'd01248408;
                12'd2299: logsin <= 24'd01249198;
                12'd2300: logsin <= 24'd01249987;
                12'd2301: logsin <= 24'd01250776;
                12'd2302: logsin <= 24'd01251565;
                12'd2303: logsin <= 24'd01252354;
                12'd2304: logsin <= 24'd01253143;
                12'd2305: logsin <= 24'd01253932;
                12'd2306: logsin <= 24'd01254720;
                12'd2307: logsin <= 24'd01255509;
                12'd2308: logsin <= 24'd01256297;
                12'd2309: logsin <= 24'd01257085;
                12'd2310: logsin <= 24'd01257874;
                12'd2311: logsin <= 24'd01258662;
                12'd2312: logsin <= 24'd01259449;
                12'd2313: logsin <= 24'd01260237;
                12'd2314: logsin <= 24'd01261025;
                12'd2315: logsin <= 24'd01261812;
                12'd2316: logsin <= 24'd01262600;
                12'd2317: logsin <= 24'd01263387;
                12'd2318: logsin <= 24'd01264174;
                12'd2319: logsin <= 24'd01264961;
                12'd2320: logsin <= 24'd01265748;
                12'd2321: logsin <= 24'd01266535;
                12'd2322: logsin <= 24'd01267321;
                12'd2323: logsin <= 24'd01268108;
                12'd2324: logsin <= 24'd01268894;
                12'd2325: logsin <= 24'd01269680;
                12'd2326: logsin <= 24'd01270467;
                12'd2327: logsin <= 24'd01271253;
                12'd2328: logsin <= 24'd01272038;
                12'd2329: logsin <= 24'd01272824;
                12'd2330: logsin <= 24'd01273610;
                12'd2331: logsin <= 24'd01274395;
                12'd2332: logsin <= 24'd01275180;
                12'd2333: logsin <= 24'd01275966;
                12'd2334: logsin <= 24'd01276751;
                12'd2335: logsin <= 24'd01277536;
                12'd2336: logsin <= 24'd01278320;
                12'd2337: logsin <= 24'd01279105;
                12'd2338: logsin <= 24'd01279889;
                12'd2339: logsin <= 24'd01280674;
                12'd2340: logsin <= 24'd01281458;
                12'd2341: logsin <= 24'd01282242;
                12'd2342: logsin <= 24'd01283026;
                12'd2343: logsin <= 24'd01283810;
                12'd2344: logsin <= 24'd01284594;
                12'd2345: logsin <= 24'd01285377;
                12'd2346: logsin <= 24'd01286161;
                12'd2347: logsin <= 24'd01286944;
                12'd2348: logsin <= 24'd01287727;
                12'd2349: logsin <= 24'd01288510;
                12'd2350: logsin <= 24'd01289293;
                12'd2351: logsin <= 24'd01290075;
                12'd2352: logsin <= 24'd01290858;
                12'd2353: logsin <= 24'd01291640;
                12'd2354: logsin <= 24'd01292423;
                12'd2355: logsin <= 24'd01293205;
                12'd2356: logsin <= 24'd01293987;
                12'd2357: logsin <= 24'd01294769;
                12'd2358: logsin <= 24'd01295550;
                12'd2359: logsin <= 24'd01296332;
                12'd2360: logsin <= 24'd01297113;
                12'd2361: logsin <= 24'd01297895;
                12'd2362: logsin <= 24'd01298676;
                12'd2363: logsin <= 24'd01299457;
                12'd2364: logsin <= 24'd01300237;
                12'd2365: logsin <= 24'd01301018;
                12'd2366: logsin <= 24'd01301799;
                12'd2367: logsin <= 24'd01302579;
                12'd2368: logsin <= 24'd01303359;
                12'd2369: logsin <= 24'd01304139;
                12'd2370: logsin <= 24'd01304919;
                12'd2371: logsin <= 24'd01305699;
                12'd2372: logsin <= 24'd01306479;
                12'd2373: logsin <= 24'd01307258;
                12'd2374: logsin <= 24'd01308037;
                12'd2375: logsin <= 24'd01308817;
                12'd2376: logsin <= 24'd01309596;
                12'd2377: logsin <= 24'd01310374;
                12'd2378: logsin <= 24'd01311153;
                12'd2379: logsin <= 24'd01311932;
                12'd2380: logsin <= 24'd01312710;
                12'd2381: logsin <= 24'd01313488;
                12'd2382: logsin <= 24'd01314266;
                12'd2383: logsin <= 24'd01315044;
                12'd2384: logsin <= 24'd01315822;
                12'd2385: logsin <= 24'd01316600;
                12'd2386: logsin <= 24'd01317377;
                12'd2387: logsin <= 24'd01318154;
                12'd2388: logsin <= 24'd01318932;
                12'd2389: logsin <= 24'd01319708;
                12'd2390: logsin <= 24'd01320485;
                12'd2391: logsin <= 24'd01321262;
                12'd2392: logsin <= 24'd01322038;
                12'd2393: logsin <= 24'd01322815;
                12'd2394: logsin <= 24'd01323591;
                12'd2395: logsin <= 24'd01324367;
                12'd2396: logsin <= 24'd01325143;
                12'd2397: logsin <= 24'd01325919;
                12'd2398: logsin <= 24'd01326694;
                12'd2399: logsin <= 24'd01327469;
                12'd2400: logsin <= 24'd01328245;
                12'd2401: logsin <= 24'd01329020;
                12'd2402: logsin <= 24'd01329794;
                12'd2403: logsin <= 24'd01330569;
                12'd2404: logsin <= 24'd01331344;
                12'd2405: logsin <= 24'd01332118;
                12'd2406: logsin <= 24'd01332892;
                12'd2407: logsin <= 24'd01333666;
                12'd2408: logsin <= 24'd01334440;
                12'd2409: logsin <= 24'd01335214;
                12'd2410: logsin <= 24'd01335987;
                12'd2411: logsin <= 24'd01336761;
                12'd2412: logsin <= 24'd01337534;
                12'd2413: logsin <= 24'd01338307;
                12'd2414: logsin <= 24'd01339080;
                12'd2415: logsin <= 24'd01339853;
                12'd2416: logsin <= 24'd01340625;
                12'd2417: logsin <= 24'd01341397;
                12'd2418: logsin <= 24'd01342170;
                12'd2419: logsin <= 24'd01342942;
                12'd2420: logsin <= 24'd01343713;
                12'd2421: logsin <= 24'd01344485;
                12'd2422: logsin <= 24'd01345256;
                12'd2423: logsin <= 24'd01346028;
                12'd2424: logsin <= 24'd01346799;
                12'd2425: logsin <= 24'd01347570;
                12'd2426: logsin <= 24'd01348341;
                12'd2427: logsin <= 24'd01349111;
                12'd2428: logsin <= 24'd01349882;
                12'd2429: logsin <= 24'd01350652;
                12'd2430: logsin <= 24'd01351422;
                12'd2431: logsin <= 24'd01352192;
                12'd2432: logsin <= 24'd01352962;
                12'd2433: logsin <= 24'd01353731;
                12'd2434: logsin <= 24'd01354500;
                12'd2435: logsin <= 24'd01355270;
                12'd2436: logsin <= 24'd01356039;
                12'd2437: logsin <= 24'd01356807;
                12'd2438: logsin <= 24'd01357576;
                12'd2439: logsin <= 24'd01358344;
                12'd2440: logsin <= 24'd01359113;
                12'd2441: logsin <= 24'd01359881;
                12'd2442: logsin <= 24'd01360649;
                12'd2443: logsin <= 24'd01361416;
                12'd2444: logsin <= 24'd01362184;
                12'd2445: logsin <= 24'd01362951;
                12'd2446: logsin <= 24'd01363718;
                12'd2447: logsin <= 24'd01364485;
                12'd2448: logsin <= 24'd01365252;
                12'd2449: logsin <= 24'd01366019;
                12'd2450: logsin <= 24'd01366785;
                12'd2451: logsin <= 24'd01367551;
                12'd2452: logsin <= 24'd01368317;
                12'd2453: logsin <= 24'd01369083;
                12'd2454: logsin <= 24'd01369849;
                12'd2455: logsin <= 24'd01370614;
                12'd2456: logsin <= 24'd01371380;
                12'd2457: logsin <= 24'd01372145;
                12'd2458: logsin <= 24'd01372910;
                12'd2459: logsin <= 24'd01373674;
                12'd2460: logsin <= 24'd01374439;
                12'd2461: logsin <= 24'd01375203;
                12'd2462: logsin <= 24'd01375967;
                12'd2463: logsin <= 24'd01376731;
                12'd2464: logsin <= 24'd01377495;
                12'd2465: logsin <= 24'd01378259;
                12'd2466: logsin <= 24'd01379022;
                12'd2467: logsin <= 24'd01379785;
                12'd2468: logsin <= 24'd01380548;
                12'd2469: logsin <= 24'd01381311;
                12'd2470: logsin <= 24'd01382074;
                12'd2471: logsin <= 24'd01382836;
                12'd2472: logsin <= 24'd01383598;
                12'd2473: logsin <= 24'd01384360;
                12'd2474: logsin <= 24'd01385122;
                12'd2475: logsin <= 24'd01385884;
                12'd2476: logsin <= 24'd01386645;
                12'd2477: logsin <= 24'd01387406;
                12'd2478: logsin <= 24'd01388167;
                12'd2479: logsin <= 24'd01388928;
                12'd2480: logsin <= 24'd01389689;
                12'd2481: logsin <= 24'd01390449;
                12'd2482: logsin <= 24'd01391209;
                12'd2483: logsin <= 24'd01391969;
                12'd2484: logsin <= 24'd01392729;
                12'd2485: logsin <= 24'd01393489;
                12'd2486: logsin <= 24'd01394248;
                12'd2487: logsin <= 24'd01395007;
                12'd2488: logsin <= 24'd01395766;
                12'd2489: logsin <= 24'd01396525;
                12'd2490: logsin <= 24'd01397283;
                12'd2491: logsin <= 24'd01398042;
                12'd2492: logsin <= 24'd01398800;
                12'd2493: logsin <= 24'd01399558;
                12'd2494: logsin <= 24'd01400316;
                12'd2495: logsin <= 24'd01401073;
                12'd2496: logsin <= 24'd01401831;
                12'd2497: logsin <= 24'd01402588;
                12'd2498: logsin <= 24'd01403345;
                12'd2499: logsin <= 24'd01404101;
                12'd2500: logsin <= 24'd01404858;
                12'd2501: logsin <= 24'd01405614;
                12'd2502: logsin <= 24'd01406370;
                12'd2503: logsin <= 24'd01407126;
                12'd2504: logsin <= 24'd01407882;
                12'd2505: logsin <= 24'd01408637;
                12'd2506: logsin <= 24'd01409392;
                12'd2507: logsin <= 24'd01410148;
                12'd2508: logsin <= 24'd01410902;
                12'd2509: logsin <= 24'd01411657;
                12'd2510: logsin <= 24'd01412411;
                12'd2511: logsin <= 24'd01413166;
                12'd2512: logsin <= 24'd01413919;
                12'd2513: logsin <= 24'd01414673;
                12'd2514: logsin <= 24'd01415427;
                12'd2515: logsin <= 24'd01416180;
                12'd2516: logsin <= 24'd01416933;
                12'd2517: logsin <= 24'd01417686;
                12'd2518: logsin <= 24'd01418439;
                12'd2519: logsin <= 24'd01419191;
                12'd2520: logsin <= 24'd01419943;
                12'd2521: logsin <= 24'd01420695;
                12'd2522: logsin <= 24'd01421447;
                12'd2523: logsin <= 24'd01422199;
                12'd2524: logsin <= 24'd01422950;
                12'd2525: logsin <= 24'd01423701;
                12'd2526: logsin <= 24'd01424452;
                12'd2527: logsin <= 24'd01425203;
                12'd2528: logsin <= 24'd01425953;
                12'd2529: logsin <= 24'd01426704;
                12'd2530: logsin <= 24'd01427454;
                12'd2531: logsin <= 24'd01428203;
                12'd2532: logsin <= 24'd01428953;
                12'd2533: logsin <= 24'd01429702;
                12'd2534: logsin <= 24'd01430451;
                12'd2535: logsin <= 24'd01431200;
                12'd2536: logsin <= 24'd01431949;
                12'd2537: logsin <= 24'd01432697;
                12'd2538: logsin <= 24'd01433446;
                12'd2539: logsin <= 24'd01434194;
                12'd2540: logsin <= 24'd01434941;
                12'd2541: logsin <= 24'd01435689;
                12'd2542: logsin <= 24'd01436436;
                12'd2543: logsin <= 24'd01437183;
                12'd2544: logsin <= 24'd01437930;
                12'd2545: logsin <= 24'd01438677;
                12'd2546: logsin <= 24'd01439423;
                12'd2547: logsin <= 24'd01440170;
                12'd2548: logsin <= 24'd01440915;
                12'd2549: logsin <= 24'd01441661;
                12'd2550: logsin <= 24'd01442407;
                12'd2551: logsin <= 24'd01443152;
                12'd2552: logsin <= 24'd01443897;
                12'd2553: logsin <= 24'd01444642;
                12'd2554: logsin <= 24'd01445386;
                12'd2555: logsin <= 24'd01446131;
                12'd2556: logsin <= 24'd01446875;
                12'd2557: logsin <= 24'd01447619;
                12'd2558: logsin <= 24'd01448362;
                12'd2559: logsin <= 24'd01449106;
                12'd2560: logsin <= 24'd01449849;
                12'd2561: logsin <= 24'd01450592;
                12'd2562: logsin <= 24'd01451334;
                12'd2563: logsin <= 24'd01452077;
                12'd2564: logsin <= 24'd01452819;
                12'd2565: logsin <= 24'd01453561;
                12'd2566: logsin <= 24'd01454303;
                12'd2567: logsin <= 24'd01455044;
                12'd2568: logsin <= 24'd01455785;
                12'd2569: logsin <= 24'd01456526;
                12'd2570: logsin <= 24'd01457267;
                12'd2571: logsin <= 24'd01458008;
                12'd2572: logsin <= 24'd01458748;
                12'd2573: logsin <= 24'd01459488;
                12'd2574: logsin <= 24'd01460228;
                12'd2575: logsin <= 24'd01460967;
                12'd2576: logsin <= 24'd01461707;
                12'd2577: logsin <= 24'd01462446;
                12'd2578: logsin <= 24'd01463185;
                12'd2579: logsin <= 24'd01463923;
                12'd2580: logsin <= 24'd01464661;
                12'd2581: logsin <= 24'd01465400;
                12'd2582: logsin <= 24'd01466137;
                12'd2583: logsin <= 24'd01466875;
                12'd2584: logsin <= 24'd01467612;
                12'd2585: logsin <= 24'd01468349;
                12'd2586: logsin <= 24'd01469086;
                12'd2587: logsin <= 24'd01469823;
                12'd2588: logsin <= 24'd01470559;
                12'd2589: logsin <= 24'd01471295;
                12'd2590: logsin <= 24'd01472031;
                12'd2591: logsin <= 24'd01472767;
                12'd2592: logsin <= 24'd01473502;
                12'd2593: logsin <= 24'd01474237;
                12'd2594: logsin <= 24'd01474972;
                12'd2595: logsin <= 24'd01475707;
                12'd2596: logsin <= 24'd01476441;
                12'd2597: logsin <= 24'd01477175;
                12'd2598: logsin <= 24'd01477909;
                12'd2599: logsin <= 24'd01478643;
                12'd2600: logsin <= 24'd01479376;
                12'd2601: logsin <= 24'd01480109;
                12'd2602: logsin <= 24'd01480842;
                12'd2603: logsin <= 24'd01481575;
                12'd2604: logsin <= 24'd01482307;
                12'd2605: logsin <= 24'd01483039;
                12'd2606: logsin <= 24'd01483771;
                12'd2607: logsin <= 24'd01484503;
                12'd2608: logsin <= 24'd01485234;
                12'd2609: logsin <= 24'd01485965;
                12'd2610: logsin <= 24'd01486696;
                12'd2611: logsin <= 24'd01487426;
                12'd2612: logsin <= 24'd01488157;
                12'd2613: logsin <= 24'd01488887;
                12'd2614: logsin <= 24'd01489617;
                12'd2615: logsin <= 24'd01490346;
                12'd2616: logsin <= 24'd01491075;
                12'd2617: logsin <= 24'd01491804;
                12'd2618: logsin <= 24'd01492533;
                12'd2619: logsin <= 24'd01493262;
                12'd2620: logsin <= 24'd01493990;
                12'd2621: logsin <= 24'd01494718;
                12'd2622: logsin <= 24'd01495445;
                12'd2623: logsin <= 24'd01496173;
                12'd2624: logsin <= 24'd01496900;
                12'd2625: logsin <= 24'd01497627;
                12'd2626: logsin <= 24'd01498354;
                12'd2627: logsin <= 24'd01499080;
                12'd2628: logsin <= 24'd01499806;
                12'd2629: logsin <= 24'd01500532;
                12'd2630: logsin <= 24'd01501257;
                12'd2631: logsin <= 24'd01501983;
                12'd2632: logsin <= 24'd01502708;
                12'd2633: logsin <= 24'd01503433;
                12'd2634: logsin <= 24'd01504157;
                12'd2635: logsin <= 24'd01504881;
                12'd2636: logsin <= 24'd01505605;
                12'd2637: logsin <= 24'd01506329;
                12'd2638: logsin <= 24'd01507052;
                12'd2639: logsin <= 24'd01507776;
                12'd2640: logsin <= 24'd01508498;
                12'd2641: logsin <= 24'd01509221;
                12'd2642: logsin <= 24'd01509943;
                12'd2643: logsin <= 24'd01510666;
                12'd2644: logsin <= 24'd01511387;
                12'd2645: logsin <= 24'd01512109;
                12'd2646: logsin <= 24'd01512830;
                12'd2647: logsin <= 24'd01513551;
                12'd2648: logsin <= 24'd01514272;
                12'd2649: logsin <= 24'd01514992;
                12'd2650: logsin <= 24'd01515712;
                12'd2651: logsin <= 24'd01516432;
                12'd2652: logsin <= 24'd01517152;
                12'd2653: logsin <= 24'd01517871;
                12'd2654: logsin <= 24'd01518590;
                12'd2655: logsin <= 24'd01519309;
                12'd2656: logsin <= 24'd01520028;
                12'd2657: logsin <= 24'd01520746;
                12'd2658: logsin <= 24'd01521464;
                12'd2659: logsin <= 24'd01522182;
                12'd2660: logsin <= 24'd01522899;
                12'd2661: logsin <= 24'd01523616;
                12'd2662: logsin <= 24'd01524333;
                12'd2663: logsin <= 24'd01525049;
                12'd2664: logsin <= 24'd01525766;
                12'd2665: logsin <= 24'd01526482;
                12'd2666: logsin <= 24'd01527197;
                12'd2667: logsin <= 24'd01527913;
                12'd2668: logsin <= 24'd01528628;
                12'd2669: logsin <= 24'd01529343;
                12'd2670: logsin <= 24'd01530058;
                12'd2671: logsin <= 24'd01530772;
                12'd2672: logsin <= 24'd01531486;
                12'd2673: logsin <= 24'd01532200;
                12'd2674: logsin <= 24'd01532913;
                12'd2675: logsin <= 24'd01533626;
                12'd2676: logsin <= 24'd01534339;
                12'd2677: logsin <= 24'd01535052;
                12'd2678: logsin <= 24'd01535764;
                12'd2679: logsin <= 24'd01536476;
                12'd2680: logsin <= 24'd01537188;
                12'd2681: logsin <= 24'd01537899;
                12'd2682: logsin <= 24'd01538610;
                12'd2683: logsin <= 24'd01539321;
                12'd2684: logsin <= 24'd01540032;
                12'd2685: logsin <= 24'd01540742;
                12'd2686: logsin <= 24'd01541452;
                12'd2687: logsin <= 24'd01542162;
                12'd2688: logsin <= 24'd01542871;
                12'd2689: logsin <= 24'd01543580;
                12'd2690: logsin <= 24'd01544289;
                12'd2691: logsin <= 24'd01544998;
                12'd2692: logsin <= 24'd01545706;
                12'd2693: logsin <= 24'd01546414;
                12'd2694: logsin <= 24'd01547122;
                12'd2695: logsin <= 24'd01547829;
                12'd2696: logsin <= 24'd01548536;
                12'd2697: logsin <= 24'd01549243;
                12'd2698: logsin <= 24'd01549950;
                12'd2699: logsin <= 24'd01550656;
                12'd2700: logsin <= 24'd01551362;
                12'd2701: logsin <= 24'd01552067;
                12'd2702: logsin <= 24'd01552773;
                12'd2703: logsin <= 24'd01553478;
                12'd2704: logsin <= 24'd01554182;
                12'd2705: logsin <= 24'd01554887;
                12'd2706: logsin <= 24'd01555591;
                12'd2707: logsin <= 24'd01556295;
                12'd2708: logsin <= 24'd01556998;
                12'd2709: logsin <= 24'd01557701;
                12'd2710: logsin <= 24'd01558404;
                12'd2711: logsin <= 24'd01559107;
                12'd2712: logsin <= 24'd01559809;
                12'd2713: logsin <= 24'd01560511;
                12'd2714: logsin <= 24'd01561213;
                12'd2715: logsin <= 24'd01561915;
                12'd2716: logsin <= 24'd01562616;
                12'd2717: logsin <= 24'd01563317;
                12'd2718: logsin <= 24'd01564017;
                12'd2719: logsin <= 24'd01564717;
                12'd2720: logsin <= 24'd01565417;
                12'd2721: logsin <= 24'd01566117;
                12'd2722: logsin <= 24'd01566816;
                12'd2723: logsin <= 24'd01567515;
                12'd2724: logsin <= 24'd01568214;
                12'd2725: logsin <= 24'd01568912;
                12'd2726: logsin <= 24'd01569610;
                12'd2727: logsin <= 24'd01570308;
                12'd2728: logsin <= 24'd01571006;
                12'd2729: logsin <= 24'd01571703;
                12'd2730: logsin <= 24'd01572400;
                12'd2731: logsin <= 24'd01573096;
                12'd2732: logsin <= 24'd01573792;
                12'd2733: logsin <= 24'd01574488;
                12'd2734: logsin <= 24'd01575184;
                12'd2735: logsin <= 24'd01575879;
                12'd2736: logsin <= 24'd01576574;
                12'd2737: logsin <= 24'd01577269;
                12'd2738: logsin <= 24'd01577963;
                12'd2739: logsin <= 24'd01578657;
                12'd2740: logsin <= 24'd01579351;
                12'd2741: logsin <= 24'd01580045;
                12'd2742: logsin <= 24'd01580738;
                12'd2743: logsin <= 24'd01581431;
                12'd2744: logsin <= 24'd01582123;
                12'd2745: logsin <= 24'd01582815;
                12'd2746: logsin <= 24'd01583507;
                12'd2747: logsin <= 24'd01584199;
                12'd2748: logsin <= 24'd01584890;
                12'd2749: logsin <= 24'd01585581;
                12'd2750: logsin <= 24'd01586272;
                12'd2751: logsin <= 24'd01586962;
                12'd2752: logsin <= 24'd01587652;
                12'd2753: logsin <= 24'd01588341;
                12'd2754: logsin <= 24'd01589031;
                12'd2755: logsin <= 24'd01589720;
                12'd2756: logsin <= 24'd01590409;
                12'd2757: logsin <= 24'd01591097;
                12'd2758: logsin <= 24'd01591785;
                12'd2759: logsin <= 24'd01592473;
                12'd2760: logsin <= 24'd01593160;
                12'd2761: logsin <= 24'd01593847;
                12'd2762: logsin <= 24'd01594534;
                12'd2763: logsin <= 24'd01595221;
                12'd2764: logsin <= 24'd01595907;
                12'd2765: logsin <= 24'd01596593;
                12'd2766: logsin <= 24'd01597278;
                12'd2767: logsin <= 24'd01597963;
                12'd2768: logsin <= 24'd01598648;
                12'd2769: logsin <= 24'd01599333;
                12'd2770: logsin <= 24'd01600017;
                12'd2771: logsin <= 24'd01600701;
                12'd2772: logsin <= 24'd01601384;
                12'd2773: logsin <= 24'd01602068;
                12'd2774: logsin <= 24'd01602751;
                12'd2775: logsin <= 24'd01603433;
                12'd2776: logsin <= 24'd01604115;
                12'd2777: logsin <= 24'd01604797;
                12'd2778: logsin <= 24'd01605479;
                12'd2779: logsin <= 24'd01606160;
                12'd2780: logsin <= 24'd01606841;
                12'd2781: logsin <= 24'd01607522;
                12'd2782: logsin <= 24'd01608202;
                12'd2783: logsin <= 24'd01608882;
                12'd2784: logsin <= 24'd01609562;
                12'd2785: logsin <= 24'd01610241;
                12'd2786: logsin <= 24'd01610920;
                12'd2787: logsin <= 24'd01611599;
                12'd2788: logsin <= 24'd01612277;
                12'd2789: logsin <= 24'd01612955;
                12'd2790: logsin <= 24'd01613633;
                12'd2791: logsin <= 24'd01614310;
                12'd2792: logsin <= 24'd01614987;
                12'd2793: logsin <= 24'd01615663;
                12'd2794: logsin <= 24'd01616340;
                12'd2795: logsin <= 24'd01617016;
                12'd2796: logsin <= 24'd01617691;
                12'd2797: logsin <= 24'd01618367;
                12'd2798: logsin <= 24'd01619042;
                12'd2799: logsin <= 24'd01619716;
                12'd2800: logsin <= 24'd01620391;
                12'd2801: logsin <= 24'd01621065;
                12'd2802: logsin <= 24'd01621738;
                12'd2803: logsin <= 24'd01622412;
                12'd2804: logsin <= 24'd01623085;
                12'd2805: logsin <= 24'd01623757;
                12'd2806: logsin <= 24'd01624429;
                12'd2807: logsin <= 24'd01625101;
                12'd2808: logsin <= 24'd01625773;
                12'd2809: logsin <= 24'd01626444;
                12'd2810: logsin <= 24'd01627115;
                12'd2811: logsin <= 24'd01627786;
                12'd2812: logsin <= 24'd01628456;
                12'd2813: logsin <= 24'd01629126;
                12'd2814: logsin <= 24'd01629796;
                12'd2815: logsin <= 24'd01630465;
                12'd2816: logsin <= 24'd01631134;
                12'd2817: logsin <= 24'd01631802;
                12'd2818: logsin <= 24'd01632470;
                12'd2819: logsin <= 24'd01633138;
                12'd2820: logsin <= 24'd01633806;
                12'd2821: logsin <= 24'd01634473;
                12'd2822: logsin <= 24'd01635140;
                12'd2823: logsin <= 24'd01635806;
                12'd2824: logsin <= 24'd01636472;
                12'd2825: logsin <= 24'd01637138;
                12'd2826: logsin <= 24'd01637803;
                12'd2827: logsin <= 24'd01638469;
                12'd2828: logsin <= 24'd01639133;
                12'd2829: logsin <= 24'd01639798;
                12'd2830: logsin <= 24'd01640462;
                12'd2831: logsin <= 24'd01641125;
                12'd2832: logsin <= 24'd01641789;
                12'd2833: logsin <= 24'd01642452;
                12'd2834: logsin <= 24'd01643114;
                12'd2835: logsin <= 24'd01643777;
                12'd2836: logsin <= 24'd01644439;
                12'd2837: logsin <= 24'd01645100;
                12'd2838: logsin <= 24'd01645762;
                12'd2839: logsin <= 24'd01646422;
                12'd2840: logsin <= 24'd01647083;
                12'd2841: logsin <= 24'd01647743;
                12'd2842: logsin <= 24'd01648403;
                12'd2843: logsin <= 24'd01649063;
                12'd2844: logsin <= 24'd01649722;
                12'd2845: logsin <= 24'd01650380;
                12'd2846: logsin <= 24'd01651039;
                12'd2847: logsin <= 24'd01651697;
                12'd2848: logsin <= 24'd01652355;
                12'd2849: logsin <= 24'd01653012;
                12'd2850: logsin <= 24'd01653669;
                12'd2851: logsin <= 24'd01654326;
                12'd2852: logsin <= 24'd01654982;
                12'd2853: logsin <= 24'd01655638;
                12'd2854: logsin <= 24'd01656293;
                12'd2855: logsin <= 24'd01656949;
                12'd2856: logsin <= 24'd01657604;
                12'd2857: logsin <= 24'd01658258;
                12'd2858: logsin <= 24'd01658912;
                12'd2859: logsin <= 24'd01659566;
                12'd2860: logsin <= 24'd01660219;
                12'd2861: logsin <= 24'd01660873;
                12'd2862: logsin <= 24'd01661525;
                12'd2863: logsin <= 24'd01662178;
                12'd2864: logsin <= 24'd01662830;
                12'd2865: logsin <= 24'd01663481;
                12'd2866: logsin <= 24'd01664132;
                12'd2867: logsin <= 24'd01664783;
                12'd2868: logsin <= 24'd01665434;
                12'd2869: logsin <= 24'd01666084;
                12'd2870: logsin <= 24'd01666734;
                12'd2871: logsin <= 24'd01667383;
                12'd2872: logsin <= 24'd01668032;
                12'd2873: logsin <= 24'd01668681;
                12'd2874: logsin <= 24'd01669330;
                12'd2875: logsin <= 24'd01669978;
                12'd2876: logsin <= 24'd01670625;
                12'd2877: logsin <= 24'd01671272;
                12'd2878: logsin <= 24'd01671919;
                12'd2879: logsin <= 24'd01672566;
                12'd2880: logsin <= 24'd01673212;
                12'd2881: logsin <= 24'd01673858;
                12'd2882: logsin <= 24'd01674503;
                12'd2883: logsin <= 24'd01675148;
                12'd2884: logsin <= 24'd01675793;
                12'd2885: logsin <= 24'd01676437;
                12'd2886: logsin <= 24'd01677081;
                12'd2887: logsin <= 24'd01677725;
                12'd2888: logsin <= 24'd01678368;
                12'd2889: logsin <= 24'd01679011;
                12'd2890: logsin <= 24'd01679653;
                12'd2891: logsin <= 24'd01680295;
                12'd2892: logsin <= 24'd01680937;
                12'd2893: logsin <= 24'd01681579;
                12'd2894: logsin <= 24'd01682219;
                12'd2895: logsin <= 24'd01682860;
                12'd2896: logsin <= 24'd01683500;
                12'd2897: logsin <= 24'd01684140;
                12'd2898: logsin <= 24'd01684780;
                12'd2899: logsin <= 24'd01685419;
                12'd2900: logsin <= 24'd01686058;
                12'd2901: logsin <= 24'd01686696;
                12'd2902: logsin <= 24'd01687334;
                12'd2903: logsin <= 24'd01687972;
                12'd2904: logsin <= 24'd01688609;
                12'd2905: logsin <= 24'd01689246;
                12'd2906: logsin <= 24'd01689882;
                12'd2907: logsin <= 24'd01690518;
                12'd2908: logsin <= 24'd01691154;
                12'd2909: logsin <= 24'd01691789;
                12'd2910: logsin <= 24'd01692424;
                12'd2911: logsin <= 24'd01693059;
                12'd2912: logsin <= 24'd01693693;
                12'd2913: logsin <= 24'd01694327;
                12'd2914: logsin <= 24'd01694960;
                12'd2915: logsin <= 24'd01695593;
                12'd2916: logsin <= 24'd01696226;
                12'd2917: logsin <= 24'd01696858;
                12'd2918: logsin <= 24'd01697490;
                12'd2919: logsin <= 24'd01698122;
                12'd2920: logsin <= 24'd01698753;
                12'd2921: logsin <= 24'd01699384;
                12'd2922: logsin <= 24'd01700014;
                12'd2923: logsin <= 24'd01700644;
                12'd2924: logsin <= 24'd01701274;
                12'd2925: logsin <= 24'd01701903;
                12'd2926: logsin <= 24'd01702532;
                12'd2927: logsin <= 24'd01703161;
                12'd2928: logsin <= 24'd01703789;
                12'd2929: logsin <= 24'd01704416;
                12'd2930: logsin <= 24'd01705044;
                12'd2931: logsin <= 24'd01705671;
                12'd2932: logsin <= 24'd01706297;
                12'd2933: logsin <= 24'd01706923;
                12'd2934: logsin <= 24'd01707549;
                12'd2935: logsin <= 24'd01708175;
                12'd2936: logsin <= 24'd01708800;
                12'd2937: logsin <= 24'd01709424;
                12'd2938: logsin <= 24'd01710048;
                12'd2939: logsin <= 24'd01710672;
                12'd2940: logsin <= 24'd01711296;
                12'd2941: logsin <= 24'd01711919;
                12'd2942: logsin <= 24'd01712541;
                12'd2943: logsin <= 24'd01713164;
                12'd2944: logsin <= 24'd01713786;
                12'd2945: logsin <= 24'd01714407;
                12'd2946: logsin <= 24'd01715028;
                12'd2947: logsin <= 24'd01715649;
                12'd2948: logsin <= 24'd01716269;
                12'd2949: logsin <= 24'd01716889;
                12'd2950: logsin <= 24'd01717509;
                12'd2951: logsin <= 24'd01718128;
                12'd2952: logsin <= 24'd01718747;
                12'd2953: logsin <= 24'd01719365;
                12'd2954: logsin <= 24'd01719983;
                12'd2955: logsin <= 24'd01720600;
                12'd2956: logsin <= 24'd01721218;
                12'd2957: logsin <= 24'd01721834;
                12'd2958: logsin <= 24'd01722451;
                12'd2959: logsin <= 24'd01723067;
                12'd2960: logsin <= 24'd01723682;
                12'd2961: logsin <= 24'd01724297;
                12'd2962: logsin <= 24'd01724912;
                12'd2963: logsin <= 24'd01725527;
                12'd2964: logsin <= 24'd01726141;
                12'd2965: logsin <= 24'd01726754;
                12'd2966: logsin <= 24'd01727367;
                12'd2967: logsin <= 24'd01727980;
                12'd2968: logsin <= 24'd01728593;
                12'd2969: logsin <= 24'd01729205;
                12'd2970: logsin <= 24'd01729816;
                12'd2971: logsin <= 24'd01730427;
                12'd2972: logsin <= 24'd01731038;
                12'd2973: logsin <= 24'd01731649;
                12'd2974: logsin <= 24'd01732259;
                12'd2975: logsin <= 24'd01732868;
                12'd2976: logsin <= 24'd01733477;
                12'd2977: logsin <= 24'd01734086;
                12'd2978: logsin <= 24'd01734695;
                12'd2979: logsin <= 24'd01735303;
                12'd2980: logsin <= 24'd01735910;
                12'd2981: logsin <= 24'd01736517;
                12'd2982: logsin <= 24'd01737124;
                12'd2983: logsin <= 24'd01737730;
                12'd2984: logsin <= 24'd01738336;
                12'd2985: logsin <= 24'd01738942;
                12'd2986: logsin <= 24'd01739547;
                12'd2987: logsin <= 24'd01740152;
                12'd2988: logsin <= 24'd01740756;
                12'd2989: logsin <= 24'd01741360;
                12'd2990: logsin <= 24'd01741963;
                12'd2991: logsin <= 24'd01742567;
                12'd2992: logsin <= 24'd01743169;
                12'd2993: logsin <= 24'd01743772;
                12'd2994: logsin <= 24'd01744373;
                12'd2995: logsin <= 24'd01744975;
                12'd2996: logsin <= 24'd01745576;
                12'd2997: logsin <= 24'd01746177;
                12'd2998: logsin <= 24'd01746777;
                12'd2999: logsin <= 24'd01747377;
                12'd3000: logsin <= 24'd01747976;
                12'd3001: logsin <= 24'd01748575;
                12'd3002: logsin <= 24'd01749174;
                12'd3003: logsin <= 24'd01749772;
                12'd3004: logsin <= 24'd01750370;
                12'd3005: logsin <= 24'd01750967;
                12'd3006: logsin <= 24'd01751564;
                12'd3007: logsin <= 24'd01752160;
                12'd3008: logsin <= 24'd01752757;
                12'd3009: logsin <= 24'd01753352;
                12'd3010: logsin <= 24'd01753948;
                12'd3011: logsin <= 24'd01754542;
                12'd3012: logsin <= 24'd01755137;
                12'd3013: logsin <= 24'd01755731;
                12'd3014: logsin <= 24'd01756325;
                12'd3015: logsin <= 24'd01756918;
                12'd3016: logsin <= 24'd01757511;
                12'd3017: logsin <= 24'd01758103;
                12'd3018: logsin <= 24'd01758695;
                12'd3019: logsin <= 24'd01759286;
                12'd3020: logsin <= 24'd01759878;
                12'd3021: logsin <= 24'd01760468;
                12'd3022: logsin <= 24'd01761059;
                12'd3023: logsin <= 24'd01761648;
                12'd3024: logsin <= 24'd01762238;
                12'd3025: logsin <= 24'd01762827;
                12'd3026: logsin <= 24'd01763416;
                12'd3027: logsin <= 24'd01764004;
                12'd3028: logsin <= 24'd01764591;
                12'd3029: logsin <= 24'd01765179;
                12'd3030: logsin <= 24'd01765766;
                12'd3031: logsin <= 24'd01766352;
                12'd3032: logsin <= 24'd01766938;
                12'd3033: logsin <= 24'd01767524;
                12'd3034: logsin <= 24'd01768109;
                12'd3035: logsin <= 24'd01768694;
                12'd3036: logsin <= 24'd01769278;
                12'd3037: logsin <= 24'd01769862;
                12'd3038: logsin <= 24'd01770446;
                12'd3039: logsin <= 24'd01771029;
                12'd3040: logsin <= 24'd01771612;
                12'd3041: logsin <= 24'd01772194;
                12'd3042: logsin <= 24'd01772776;
                12'd3043: logsin <= 24'd01773357;
                12'd3044: logsin <= 24'd01773938;
                12'd3045: logsin <= 24'd01774519;
                12'd3046: logsin <= 24'd01775099;
                12'd3047: logsin <= 24'd01775679;
                12'd3048: logsin <= 24'd01776258;
                12'd3049: logsin <= 24'd01776837;
                12'd3050: logsin <= 24'd01777415;
                12'd3051: logsin <= 24'd01777993;
                12'd3052: logsin <= 24'd01778571;
                12'd3053: logsin <= 24'd01779148;
                12'd3054: logsin <= 24'd01779724;
                12'd3055: logsin <= 24'd01780301;
                12'd3056: logsin <= 24'd01780877;
                12'd3057: logsin <= 24'd01781452;
                12'd3058: logsin <= 24'd01782027;
                12'd3059: logsin <= 24'd01782602;
                12'd3060: logsin <= 24'd01783176;
                12'd3061: logsin <= 24'd01783749;
                12'd3062: logsin <= 24'd01784323;
                12'd3063: logsin <= 24'd01784895;
                12'd3064: logsin <= 24'd01785468;
                12'd3065: logsin <= 24'd01786040;
                12'd3066: logsin <= 24'd01786611;
                12'd3067: logsin <= 24'd01787182;
                12'd3068: logsin <= 24'd01787753;
                12'd3069: logsin <= 24'd01788323;
                12'd3070: logsin <= 24'd01788893;
                12'd3071: logsin <= 24'd01789462;
                12'd3072: logsin <= 24'd01790031;
                12'd3073: logsin <= 24'd01790600;
                12'd3074: logsin <= 24'd01791168;
                12'd3075: logsin <= 24'd01791735;
                12'd3076: logsin <= 24'd01792302;
                12'd3077: logsin <= 24'd01792869;
                12'd3078: logsin <= 24'd01793435;
                12'd3079: logsin <= 24'd01794001;
                12'd3080: logsin <= 24'd01794567;
                12'd3081: logsin <= 24'd01795132;
                12'd3082: logsin <= 24'd01795696;
                12'd3083: logsin <= 24'd01796260;
                12'd3084: logsin <= 24'd01796824;
                12'd3085: logsin <= 24'd01797387;
                12'd3086: logsin <= 24'd01797950;
                12'd3087: logsin <= 24'd01798512;
                12'd3088: logsin <= 24'd01799074;
                12'd3089: logsin <= 24'd01799636;
                12'd3090: logsin <= 24'd01800197;
                12'd3091: logsin <= 24'd01800757;
                12'd3092: logsin <= 24'd01801317;
                12'd3093: logsin <= 24'd01801877;
                12'd3094: logsin <= 24'd01802436;
                12'd3095: logsin <= 24'd01802995;
                12'd3096: logsin <= 24'd01803553;
                12'd3097: logsin <= 24'd01804111;
                12'd3098: logsin <= 24'd01804669;
                12'd3099: logsin <= 24'd01805226;
                12'd3100: logsin <= 24'd01805782;
                12'd3101: logsin <= 24'd01806338;
                12'd3102: logsin <= 24'd01806894;
                12'd3103: logsin <= 24'd01807449;
                12'd3104: logsin <= 24'd01808004;
                12'd3105: logsin <= 24'd01808558;
                12'd3106: logsin <= 24'd01809112;
                12'd3107: logsin <= 24'd01809666;
                12'd3108: logsin <= 24'd01810219;
                12'd3109: logsin <= 24'd01810771;
                12'd3110: logsin <= 24'd01811323;
                12'd3111: logsin <= 24'd01811875;
                12'd3112: logsin <= 24'd01812426;
                12'd3113: logsin <= 24'd01812977;
                12'd3114: logsin <= 24'd01813527;
                12'd3115: logsin <= 24'd01814077;
                12'd3116: logsin <= 24'd01814627;
                12'd3117: logsin <= 24'd01815176;
                12'd3118: logsin <= 24'd01815724;
                12'd3119: logsin <= 24'd01816272;
                12'd3120: logsin <= 24'd01816820;
                12'd3121: logsin <= 24'd01817367;
                12'd3122: logsin <= 24'd01817914;
                12'd3123: logsin <= 24'd01818460;
                12'd3124: logsin <= 24'd01819006;
                12'd3125: logsin <= 24'd01819551;
                12'd3126: logsin <= 24'd01820096;
                12'd3127: logsin <= 24'd01820640;
                12'd3128: logsin <= 24'd01821184;
                12'd3129: logsin <= 24'd01821728;
                12'd3130: logsin <= 24'd01822271;
                12'd3131: logsin <= 24'd01822813;
                12'd3132: logsin <= 24'd01823356;
                12'd3133: logsin <= 24'd01823897;
                12'd3134: logsin <= 24'd01824438;
                12'd3135: logsin <= 24'd01824979;
                12'd3136: logsin <= 24'd01825520;
                12'd3137: logsin <= 24'd01826059;
                12'd3138: logsin <= 24'd01826599;
                12'd3139: logsin <= 24'd01827138;
                12'd3140: logsin <= 24'd01827676;
                12'd3141: logsin <= 24'd01828214;
                12'd3142: logsin <= 24'd01828752;
                12'd3143: logsin <= 24'd01829289;
                12'd3144: logsin <= 24'd01829826;
                12'd3145: logsin <= 24'd01830362;
                12'd3146: logsin <= 24'd01830898;
                12'd3147: logsin <= 24'd01831433;
                12'd3148: logsin <= 24'd01831968;
                12'd3149: logsin <= 24'd01832502;
                12'd3150: logsin <= 24'd01833036;
                12'd3151: logsin <= 24'd01833569;
                12'd3152: logsin <= 24'd01834102;
                12'd3153: logsin <= 24'd01834635;
                12'd3154: logsin <= 24'd01835167;
                12'd3155: logsin <= 24'd01835699;
                12'd3156: logsin <= 24'd01836230;
                12'd3157: logsin <= 24'd01836760;
                12'd3158: logsin <= 24'd01837291;
                12'd3159: logsin <= 24'd01837820;
                12'd3160: logsin <= 24'd01838350;
                12'd3161: logsin <= 24'd01838878;
                12'd3162: logsin <= 24'd01839407;
                12'd3163: logsin <= 24'd01839935;
                12'd3164: logsin <= 24'd01840462;
                12'd3165: logsin <= 24'd01840989;
                12'd3166: logsin <= 24'd01841515;
                12'd3167: logsin <= 24'd01842041;
                12'd3168: logsin <= 24'd01842567;
                12'd3169: logsin <= 24'd01843092;
                12'd3170: logsin <= 24'd01843617;
                12'd3171: logsin <= 24'd01844141;
                12'd3172: logsin <= 24'd01844665;
                12'd3173: logsin <= 24'd01845188;
                12'd3174: logsin <= 24'd01845710;
                12'd3175: logsin <= 24'd01846233;
                12'd3176: logsin <= 24'd01846755;
                12'd3177: logsin <= 24'd01847276;
                12'd3178: logsin <= 24'd01847797;
                12'd3179: logsin <= 24'd01848317;
                12'd3180: logsin <= 24'd01848837;
                12'd3181: logsin <= 24'd01849357;
                12'd3182: logsin <= 24'd01849875;
                12'd3183: logsin <= 24'd01850394;
                12'd3184: logsin <= 24'd01850912;
                12'd3185: logsin <= 24'd01851430;
                12'd3186: logsin <= 24'd01851947;
                12'd3187: logsin <= 24'd01852463;
                12'd3188: logsin <= 24'd01852979;
                12'd3189: logsin <= 24'd01853495;
                12'd3190: logsin <= 24'd01854010;
                12'd3191: logsin <= 24'd01854525;
                12'd3192: logsin <= 24'd01855039;
                12'd3193: logsin <= 24'd01855553;
                12'd3194: logsin <= 24'd01856066;
                12'd3195: logsin <= 24'd01856579;
                12'd3196: logsin <= 24'd01857092;
                12'd3197: logsin <= 24'd01857603;
                12'd3198: logsin <= 24'd01858115;
                12'd3199: logsin <= 24'd01858626;
                12'd3200: logsin <= 24'd01859136;
                12'd3201: logsin <= 24'd01859646;
                12'd3202: logsin <= 24'd01860156;
                12'd3203: logsin <= 24'd01860665;
                12'd3204: logsin <= 24'd01861173;
                12'd3205: logsin <= 24'd01861681;
                12'd3206: logsin <= 24'd01862189;
                12'd3207: logsin <= 24'd01862696;
                12'd3208: logsin <= 24'd01863203;
                12'd3209: logsin <= 24'd01863709;
                12'd3210: logsin <= 24'd01864214;
                12'd3211: logsin <= 24'd01864720;
                12'd3212: logsin <= 24'd01865224;
                12'd3213: logsin <= 24'd01865729;
                12'd3214: logsin <= 24'd01866232;
                12'd3215: logsin <= 24'd01866736;
                12'd3216: logsin <= 24'd01867238;
                12'd3217: logsin <= 24'd01867741;
                12'd3218: logsin <= 24'd01868242;
                12'd3219: logsin <= 24'd01868744;
                12'd3220: logsin <= 24'd01869245;
                12'd3221: logsin <= 24'd01869745;
                12'd3222: logsin <= 24'd01870245;
                12'd3223: logsin <= 24'd01870744;
                12'd3224: logsin <= 24'd01871243;
                12'd3225: logsin <= 24'd01871742;
                12'd3226: logsin <= 24'd01872240;
                12'd3227: logsin <= 24'd01872737;
                12'd3228: logsin <= 24'd01873234;
                12'd3229: logsin <= 24'd01873731;
                12'd3230: logsin <= 24'd01874227;
                12'd3231: logsin <= 24'd01874722;
                12'd3232: logsin <= 24'd01875217;
                12'd3233: logsin <= 24'd01875712;
                12'd3234: logsin <= 24'd01876206;
                12'd3235: logsin <= 24'd01876699;
                12'd3236: logsin <= 24'd01877192;
                12'd3237: logsin <= 24'd01877685;
                12'd3238: logsin <= 24'd01878177;
                12'd3239: logsin <= 24'd01878669;
                12'd3240: logsin <= 24'd01879160;
                12'd3241: logsin <= 24'd01879651;
                12'd3242: logsin <= 24'd01880141;
                12'd3243: logsin <= 24'd01880630;
                12'd3244: logsin <= 24'd01881120;
                12'd3245: logsin <= 24'd01881608;
                12'd3246: logsin <= 24'd01882097;
                12'd3247: logsin <= 24'd01882584;
                12'd3248: logsin <= 24'd01883071;
                12'd3249: logsin <= 24'd01883558;
                12'd3250: logsin <= 24'd01884044;
                12'd3251: logsin <= 24'd01884530;
                12'd3252: logsin <= 24'd01885015;
                12'd3253: logsin <= 24'd01885500;
                12'd3254: logsin <= 24'd01885985;
                12'd3255: logsin <= 24'd01886468;
                12'd3256: logsin <= 24'd01886952;
                12'd3257: logsin <= 24'd01887434;
                12'd3258: logsin <= 24'd01887917;
                12'd3259: logsin <= 24'd01888399;
                12'd3260: logsin <= 24'd01888880;
                12'd3261: logsin <= 24'd01889361;
                12'd3262: logsin <= 24'd01889841;
                12'd3263: logsin <= 24'd01890321;
                12'd3264: logsin <= 24'd01890800;
                12'd3265: logsin <= 24'd01891279;
                12'd3266: logsin <= 24'd01891757;
                12'd3267: logsin <= 24'd01892235;
                12'd3268: logsin <= 24'd01892713;
                12'd3269: logsin <= 24'd01893189;
                12'd3270: logsin <= 24'd01893666;
                12'd3271: logsin <= 24'd01894142;
                12'd3272: logsin <= 24'd01894617;
                12'd3273: logsin <= 24'd01895092;
                12'd3274: logsin <= 24'd01895566;
                12'd3275: logsin <= 24'd01896040;
                12'd3276: logsin <= 24'd01896513;
                12'd3277: logsin <= 24'd01896986;
                12'd3278: logsin <= 24'd01897459;
                12'd3279: logsin <= 24'd01897931;
                12'd3280: logsin <= 24'd01898402;
                12'd3281: logsin <= 24'd01898873;
                12'd3282: logsin <= 24'd01899343;
                12'd3283: logsin <= 24'd01899813;
                12'd3284: logsin <= 24'd01900282;
                12'd3285: logsin <= 24'd01900751;
                12'd3286: logsin <= 24'd01901220;
                12'd3287: logsin <= 24'd01901688;
                12'd3288: logsin <= 24'd01902155;
                12'd3289: logsin <= 24'd01902622;
                12'd3290: logsin <= 24'd01903088;
                12'd3291: logsin <= 24'd01903554;
                12'd3292: logsin <= 24'd01904019;
                12'd3293: logsin <= 24'd01904484;
                12'd3294: logsin <= 24'd01904949;
                12'd3295: logsin <= 24'd01905412;
                12'd3296: logsin <= 24'd01905876;
                12'd3297: logsin <= 24'd01906339;
                12'd3298: logsin <= 24'd01906801;
                12'd3299: logsin <= 24'd01907263;
                12'd3300: logsin <= 24'd01907724;
                12'd3301: logsin <= 24'd01908185;
                12'd3302: logsin <= 24'd01908645;
                12'd3303: logsin <= 24'd01909105;
                12'd3304: logsin <= 24'd01909564;
                12'd3305: logsin <= 24'd01910023;
                12'd3306: logsin <= 24'd01910481;
                12'd3307: logsin <= 24'd01910939;
                12'd3308: logsin <= 24'd01911397;
                12'd3309: logsin <= 24'd01911853;
                12'd3310: logsin <= 24'd01912310;
                12'd3311: logsin <= 24'd01912765;
                12'd3312: logsin <= 24'd01913221;
                12'd3313: logsin <= 24'd01913675;
                12'd3314: logsin <= 24'd01914130;
                12'd3315: logsin <= 24'd01914583;
                12'd3316: logsin <= 24'd01915036;
                12'd3317: logsin <= 24'd01915489;
                12'd3318: logsin <= 24'd01915941;
                12'd3319: logsin <= 24'd01916393;
                12'd3320: logsin <= 24'd01916844;
                12'd3321: logsin <= 24'd01917295;
                12'd3322: logsin <= 24'd01917745;
                12'd3323: logsin <= 24'd01918195;
                12'd3324: logsin <= 24'd01918644;
                12'd3325: logsin <= 24'd01919092;
                12'd3326: logsin <= 24'd01919540;
                12'd3327: logsin <= 24'd01919988;
                12'd3328: logsin <= 24'd01920435;
                12'd3329: logsin <= 24'd01920882;
                12'd3330: logsin <= 24'd01921328;
                12'd3331: logsin <= 24'd01921773;
                12'd3332: logsin <= 24'd01922218;
                12'd3333: logsin <= 24'd01922663;
                12'd3334: logsin <= 24'd01923107;
                12'd3335: logsin <= 24'd01923550;
                12'd3336: logsin <= 24'd01923993;
                12'd3337: logsin <= 24'd01924436;
                12'd3338: logsin <= 24'd01924878;
                12'd3339: logsin <= 24'd01925319;
                12'd3340: logsin <= 24'd01925760;
                12'd3341: logsin <= 24'd01926200;
                12'd3342: logsin <= 24'd01926640;
                12'd3343: logsin <= 24'd01927079;
                12'd3344: logsin <= 24'd01927518;
                12'd3345: logsin <= 24'd01927957;
                12'd3346: logsin <= 24'd01928394;
                12'd3347: logsin <= 24'd01928832;
                12'd3348: logsin <= 24'd01929268;
                12'd3349: logsin <= 24'd01929705;
                12'd3350: logsin <= 24'd01930140;
                12'd3351: logsin <= 24'd01930576;
                12'd3352: logsin <= 24'd01931010;
                12'd3353: logsin <= 24'd01931445;
                12'd3354: logsin <= 24'd01931878;
                12'd3355: logsin <= 24'd01932311;
                12'd3356: logsin <= 24'd01932744;
                12'd3357: logsin <= 24'd01933176;
                12'd3358: logsin <= 24'd01933608;
                12'd3359: logsin <= 24'd01934039;
                12'd3360: logsin <= 24'd01934469;
                12'd3361: logsin <= 24'd01934899;
                12'd3362: logsin <= 24'd01935329;
                12'd3363: logsin <= 24'd01935758;
                12'd3364: logsin <= 24'd01936186;
                12'd3365: logsin <= 24'd01936614;
                12'd3366: logsin <= 24'd01937041;
                12'd3367: logsin <= 24'd01937468;
                12'd3368: logsin <= 24'd01937895;
                12'd3369: logsin <= 24'd01938320;
                12'd3370: logsin <= 24'd01938746;
                12'd3371: logsin <= 24'd01939171;
                12'd3372: logsin <= 24'd01939595;
                12'd3373: logsin <= 24'd01940019;
                12'd3374: logsin <= 24'd01940442;
                12'd3375: logsin <= 24'd01940864;
                12'd3376: logsin <= 24'd01941287;
                12'd3377: logsin <= 24'd01941708;
                12'd3378: logsin <= 24'd01942129;
                12'd3379: logsin <= 24'd01942550;
                12'd3380: logsin <= 24'd01942970;
                12'd3381: logsin <= 24'd01943390;
                12'd3382: logsin <= 24'd01943809;
                12'd3383: logsin <= 24'd01944227;
                12'd3384: logsin <= 24'd01944645;
                12'd3385: logsin <= 24'd01945062;
                12'd3386: logsin <= 24'd01945479;
                12'd3387: logsin <= 24'd01945896;
                12'd3388: logsin <= 24'd01946312;
                12'd3389: logsin <= 24'd01946727;
                12'd3390: logsin <= 24'd01947142;
                12'd3391: logsin <= 24'd01947556;
                12'd3392: logsin <= 24'd01947970;
                12'd3393: logsin <= 24'd01948383;
                12'd3394: logsin <= 24'd01948796;
                12'd3395: logsin <= 24'd01949208;
                12'd3396: logsin <= 24'd01949619;
                12'd3397: logsin <= 24'd01950030;
                12'd3398: logsin <= 24'd01950441;
                12'd3399: logsin <= 24'd01950851;
                12'd3400: logsin <= 24'd01951260;
                12'd3401: logsin <= 24'd01951669;
                12'd3402: logsin <= 24'd01952078;
                12'd3403: logsin <= 24'd01952486;
                12'd3404: logsin <= 24'd01952893;
                12'd3405: logsin <= 24'd01953300;
                12'd3406: logsin <= 24'd01953706;
                12'd3407: logsin <= 24'd01954112;
                12'd3408: logsin <= 24'd01954517;
                12'd3409: logsin <= 24'd01954922;
                12'd3410: logsin <= 24'd01955326;
                12'd3411: logsin <= 24'd01955730;
                12'd3412: logsin <= 24'd01956133;
                12'd3413: logsin <= 24'd01956535;
                12'd3414: logsin <= 24'd01956937;
                12'd3415: logsin <= 24'd01957339;
                12'd3416: logsin <= 24'd01957740;
                12'd3417: logsin <= 24'd01958140;
                12'd3418: logsin <= 24'd01958540;
                12'd3419: logsin <= 24'd01958940;
                12'd3420: logsin <= 24'd01959338;
                12'd3421: logsin <= 24'd01959737;
                12'd3422: logsin <= 24'd01960134;
                12'd3423: logsin <= 24'd01960532;
                12'd3424: logsin <= 24'd01960928;
                12'd3425: logsin <= 24'd01961324;
                12'd3426: logsin <= 24'd01961720;
                12'd3427: logsin <= 24'd01962115;
                12'd3428: logsin <= 24'd01962510;
                12'd3429: logsin <= 24'd01962904;
                12'd3430: logsin <= 24'd01963297;
                12'd3431: logsin <= 24'd01963690;
                12'd3432: logsin <= 24'd01964082;
                12'd3433: logsin <= 24'd01964474;
                12'd3434: logsin <= 24'd01964866;
                12'd3435: logsin <= 24'd01965256;
                12'd3436: logsin <= 24'd01965647;
                12'd3437: logsin <= 24'd01966036;
                12'd3438: logsin <= 24'd01966425;
                12'd3439: logsin <= 24'd01966814;
                12'd3440: logsin <= 24'd01967202;
                12'd3441: logsin <= 24'd01967590;
                12'd3442: logsin <= 24'd01967977;
                12'd3443: logsin <= 24'd01968363;
                12'd3444: logsin <= 24'd01968749;
                12'd3445: logsin <= 24'd01969134;
                12'd3446: logsin <= 24'd01969519;
                12'd3447: logsin <= 24'd01969903;
                12'd3448: logsin <= 24'd01970287;
                12'd3449: logsin <= 24'd01970670;
                12'd3450: logsin <= 24'd01971053;
                12'd3451: logsin <= 24'd01971435;
                12'd3452: logsin <= 24'd01971817;
                12'd3453: logsin <= 24'd01972198;
                12'd3454: logsin <= 24'd01972578;
                12'd3455: logsin <= 24'd01972958;
                12'd3456: logsin <= 24'd01973337;
                12'd3457: logsin <= 24'd01973716;
                12'd3458: logsin <= 24'd01974095;
                12'd3459: logsin <= 24'd01974472;
                12'd3460: logsin <= 24'd01974850;
                12'd3461: logsin <= 24'd01975226;
                12'd3462: logsin <= 24'd01975602;
                12'd3463: logsin <= 24'd01975978;
                12'd3464: logsin <= 24'd01976353;
                12'd3465: logsin <= 24'd01976727;
                12'd3466: logsin <= 24'd01977101;
                12'd3467: logsin <= 24'd01977475;
                12'd3468: logsin <= 24'd01977848;
                12'd3469: logsin <= 24'd01978220;
                12'd3470: logsin <= 24'd01978592;
                12'd3471: logsin <= 24'd01978963;
                12'd3472: logsin <= 24'd01979334;
                12'd3473: logsin <= 24'd01979704;
                12'd3474: logsin <= 24'd01980073;
                12'd3475: logsin <= 24'd01980442;
                12'd3476: logsin <= 24'd01980811;
                12'd3477: logsin <= 24'd01981179;
                12'd3478: logsin <= 24'd01981546;
                12'd3479: logsin <= 24'd01981913;
                12'd3480: logsin <= 24'd01982279;
                12'd3481: logsin <= 24'd01982645;
                12'd3482: logsin <= 24'd01983010;
                12'd3483: logsin <= 24'd01983375;
                12'd3484: logsin <= 24'd01983739;
                12'd3485: logsin <= 24'd01984102;
                12'd3486: logsin <= 24'd01984465;
                12'd3487: logsin <= 24'd01984828;
                12'd3488: logsin <= 24'd01985190;
                12'd3489: logsin <= 24'd01985551;
                12'd3490: logsin <= 24'd01985912;
                12'd3491: logsin <= 24'd01986272;
                12'd3492: logsin <= 24'd01986632;
                12'd3493: logsin <= 24'd01986991;
                12'd3494: logsin <= 24'd01987349;
                12'd3495: logsin <= 24'd01987707;
                12'd3496: logsin <= 24'd01988065;
                12'd3497: logsin <= 24'd01988422;
                12'd3498: logsin <= 24'd01988778;
                12'd3499: logsin <= 24'd01989134;
                12'd3500: logsin <= 24'd01989489;
                12'd3501: logsin <= 24'd01989844;
                12'd3502: logsin <= 24'd01990198;
                12'd3503: logsin <= 24'd01990551;
                12'd3504: logsin <= 24'd01990904;
                12'd3505: logsin <= 24'd01991257;
                12'd3506: logsin <= 24'd01991609;
                12'd3507: logsin <= 24'd01991960;
                12'd3508: logsin <= 24'd01992311;
                12'd3509: logsin <= 24'd01992661;
                12'd3510: logsin <= 24'd01993011;
                12'd3511: logsin <= 24'd01993360;
                12'd3512: logsin <= 24'd01993709;
                12'd3513: logsin <= 24'd01994057;
                12'd3514: logsin <= 24'd01994404;
                12'd3515: logsin <= 24'd01994751;
                12'd3516: logsin <= 24'd01995098;
                12'd3517: logsin <= 24'd01995443;
                12'd3518: logsin <= 24'd01995789;
                12'd3519: logsin <= 24'd01996133;
                12'd3520: logsin <= 24'd01996477;
                12'd3521: logsin <= 24'd01996821;
                12'd3522: logsin <= 24'd01997164;
                12'd3523: logsin <= 24'd01997507;
                12'd3524: logsin <= 24'd01997848;
                12'd3525: logsin <= 24'd01998190;
                12'd3526: logsin <= 24'd01998531;
                12'd3527: logsin <= 24'd01998871;
                12'd3528: logsin <= 24'd01999210;
                12'd3529: logsin <= 24'd01999550;
                12'd3530: logsin <= 24'd01999888;
                12'd3531: logsin <= 24'd02000226;
                12'd3532: logsin <= 24'd02000564;
                12'd3533: logsin <= 24'd02000900;
                12'd3534: logsin <= 24'd02001237;
                12'd3535: logsin <= 24'd02001573;
                12'd3536: logsin <= 24'd02001908;
                12'd3537: logsin <= 24'd02002242;
                12'd3538: logsin <= 24'd02002576;
                12'd3539: logsin <= 24'd02002910;
                12'd3540: logsin <= 24'd02003243;
                12'd3541: logsin <= 24'd02003575;
                12'd3542: logsin <= 24'd02003907;
                12'd3543: logsin <= 24'd02004238;
                12'd3544: logsin <= 24'd02004569;
                12'd3545: logsin <= 24'd02004899;
                12'd3546: logsin <= 24'd02005229;
                12'd3547: logsin <= 24'd02005558;
                12'd3548: logsin <= 24'd02005886;
                12'd3549: logsin <= 24'd02006214;
                12'd3550: logsin <= 24'd02006541;
                12'd3551: logsin <= 24'd02006868;
                12'd3552: logsin <= 24'd02007194;
                12'd3553: logsin <= 24'd02007520;
                12'd3554: logsin <= 24'd02007845;
                12'd3555: logsin <= 24'd02008170;
                12'd3556: logsin <= 24'd02008494;
                12'd3557: logsin <= 24'd02008817;
                12'd3558: logsin <= 24'd02009140;
                12'd3559: logsin <= 24'd02009462;
                12'd3560: logsin <= 24'd02009784;
                12'd3561: logsin <= 24'd02010105;
                12'd3562: logsin <= 24'd02010425;
                12'd3563: logsin <= 24'd02010745;
                12'd3564: logsin <= 24'd02011065;
                12'd3565: logsin <= 24'd02011384;
                12'd3566: logsin <= 24'd02011702;
                12'd3567: logsin <= 24'd02012020;
                12'd3568: logsin <= 24'd02012337;
                12'd3569: logsin <= 24'd02012653;
                12'd3570: logsin <= 24'd02012969;
                12'd3571: logsin <= 24'd02013285;
                12'd3572: logsin <= 24'd02013600;
                12'd3573: logsin <= 24'd02013914;
                12'd3574: logsin <= 24'd02014228;
                12'd3575: logsin <= 24'd02014541;
                12'd3576: logsin <= 24'd02014854;
                12'd3577: logsin <= 24'd02015166;
                12'd3578: logsin <= 24'd02015477;
                12'd3579: logsin <= 24'd02015788;
                12'd3580: logsin <= 24'd02016098;
                12'd3581: logsin <= 24'd02016408;
                12'd3582: logsin <= 24'd02016717;
                12'd3583: logsin <= 24'd02017026;
                12'd3584: logsin <= 24'd02017334;
                12'd3585: logsin <= 24'd02017641;
                12'd3586: logsin <= 24'd02017948;
                12'd3587: logsin <= 24'd02018255;
                12'd3588: logsin <= 24'd02018560;
                12'd3589: logsin <= 24'd02018866;
                12'd3590: logsin <= 24'd02019170;
                12'd3591: logsin <= 24'd02019474;
                12'd3592: logsin <= 24'd02019778;
                12'd3593: logsin <= 24'd02020081;
                12'd3594: logsin <= 24'd02020383;
                12'd3595: logsin <= 24'd02020685;
                12'd3596: logsin <= 24'd02020986;
                12'd3597: logsin <= 24'd02021287;
                12'd3598: logsin <= 24'd02021587;
                12'd3599: logsin <= 24'd02021886;
                12'd3600: logsin <= 24'd02022185;
                12'd3601: logsin <= 24'd02022484;
                12'd3602: logsin <= 24'd02022781;
                12'd3603: logsin <= 24'd02023079;
                12'd3604: logsin <= 24'd02023375;
                12'd3605: logsin <= 24'd02023671;
                12'd3606: logsin <= 24'd02023967;
                12'd3607: logsin <= 24'd02024262;
                12'd3608: logsin <= 24'd02024556;
                12'd3609: logsin <= 24'd02024850;
                12'd3610: logsin <= 24'd02025143;
                12'd3611: logsin <= 24'd02025435;
                12'd3612: logsin <= 24'd02025727;
                12'd3613: logsin <= 24'd02026019;
                12'd3614: logsin <= 24'd02026310;
                12'd3615: logsin <= 24'd02026600;
                12'd3616: logsin <= 24'd02026890;
                12'd3617: logsin <= 24'd02027179;
                12'd3618: logsin <= 24'd02027468;
                12'd3619: logsin <= 24'd02027756;
                12'd3620: logsin <= 24'd02028043;
                12'd3621: logsin <= 24'd02028330;
                12'd3622: logsin <= 24'd02028616;
                12'd3623: logsin <= 24'd02028902;
                12'd3624: logsin <= 24'd02029187;
                12'd3625: logsin <= 24'd02029472;
                12'd3626: logsin <= 24'd02029756;
                12'd3627: logsin <= 24'd02030039;
                12'd3628: logsin <= 24'd02030322;
                12'd3629: logsin <= 24'd02030604;
                12'd3630: logsin <= 24'd02030886;
                12'd3631: logsin <= 24'd02031167;
                12'd3632: logsin <= 24'd02031447;
                12'd3633: logsin <= 24'd02031727;
                12'd3634: logsin <= 24'd02032006;
                12'd3635: logsin <= 24'd02032285;
                12'd3636: logsin <= 24'd02032563;
                12'd3637: logsin <= 24'd02032841;
                12'd3638: logsin <= 24'd02033118;
                12'd3639: logsin <= 24'd02033395;
                12'd3640: logsin <= 24'd02033670;
                12'd3641: logsin <= 24'd02033946;
                12'd3642: logsin <= 24'd02034220;
                12'd3643: logsin <= 24'd02034495;
                12'd3644: logsin <= 24'd02034768;
                12'd3645: logsin <= 24'd02035041;
                12'd3646: logsin <= 24'd02035313;
                12'd3647: logsin <= 24'd02035585;
                12'd3648: logsin <= 24'd02035857;
                12'd3649: logsin <= 24'd02036127;
                12'd3650: logsin <= 24'd02036397;
                12'd3651: logsin <= 24'd02036667;
                12'd3652: logsin <= 24'd02036936;
                12'd3653: logsin <= 24'd02037204;
                12'd3654: logsin <= 24'd02037472;
                12'd3655: logsin <= 24'd02037739;
                12'd3656: logsin <= 24'd02038005;
                12'd3657: logsin <= 24'd02038271;
                12'd3658: logsin <= 24'd02038537;
                12'd3659: logsin <= 24'd02038802;
                12'd3660: logsin <= 24'd02039066;
                12'd3661: logsin <= 24'd02039330;
                12'd3662: logsin <= 24'd02039593;
                12'd3663: logsin <= 24'd02039855;
                12'd3664: logsin <= 24'd02040117;
                12'd3665: logsin <= 24'd02040378;
                12'd3666: logsin <= 24'd02040639;
                12'd3667: logsin <= 24'd02040899;
                12'd3668: logsin <= 24'd02041159;
                12'd3669: logsin <= 24'd02041418;
                12'd3670: logsin <= 24'd02041676;
                12'd3671: logsin <= 24'd02041934;
                12'd3672: logsin <= 24'd02042192;
                12'd3673: logsin <= 24'd02042448;
                12'd3674: logsin <= 24'd02042704;
                12'd3675: logsin <= 24'd02042960;
                12'd3676: logsin <= 24'd02043215;
                12'd3677: logsin <= 24'd02043469;
                12'd3678: logsin <= 24'd02043723;
                12'd3679: logsin <= 24'd02043976;
                12'd3680: logsin <= 24'd02044228;
                12'd3681: logsin <= 24'd02044480;
                12'd3682: logsin <= 24'd02044732;
                12'd3683: logsin <= 24'd02044983;
                12'd3684: logsin <= 24'd02045233;
                12'd3685: logsin <= 24'd02045483;
                12'd3686: logsin <= 24'd02045732;
                12'd3687: logsin <= 24'd02045980;
                12'd3688: logsin <= 24'd02046228;
                12'd3689: logsin <= 24'd02046475;
                12'd3690: logsin <= 24'd02046722;
                12'd3691: logsin <= 24'd02046968;
                12'd3692: logsin <= 24'd02047214;
                12'd3693: logsin <= 24'd02047459;
                12'd3694: logsin <= 24'd02047703;
                12'd3695: logsin <= 24'd02047947;
                12'd3696: logsin <= 24'd02048190;
                12'd3697: logsin <= 24'd02048432;
                12'd3698: logsin <= 24'd02048674;
                12'd3699: logsin <= 24'd02048916;
                12'd3700: logsin <= 24'd02049157;
                12'd3701: logsin <= 24'd02049397;
                12'd3702: logsin <= 24'd02049637;
                12'd3703: logsin <= 24'd02049876;
                12'd3704: logsin <= 24'd02050114;
                12'd3705: logsin <= 24'd02050352;
                12'd3706: logsin <= 24'd02050589;
                12'd3707: logsin <= 24'd02050826;
                12'd3708: logsin <= 24'd02051062;
                12'd3709: logsin <= 24'd02051298;
                12'd3710: logsin <= 24'd02051533;
                12'd3711: logsin <= 24'd02051767;
                12'd3712: logsin <= 24'd02052001;
                12'd3713: logsin <= 24'd02052234;
                12'd3714: logsin <= 24'd02052466;
                12'd3715: logsin <= 24'd02052698;
                12'd3716: logsin <= 24'd02052930;
                12'd3717: logsin <= 24'd02053161;
                12'd3718: logsin <= 24'd02053391;
                12'd3719: logsin <= 24'd02053620;
                12'd3720: logsin <= 24'd02053849;
                12'd3721: logsin <= 24'd02054078;
                12'd3722: logsin <= 24'd02054306;
                12'd3723: logsin <= 24'd02054533;
                12'd3724: logsin <= 24'd02054760;
                12'd3725: logsin <= 24'd02054986;
                12'd3726: logsin <= 24'd02055211;
                12'd3727: logsin <= 24'd02055436;
                12'd3728: logsin <= 24'd02055660;
                12'd3729: logsin <= 24'd02055884;
                12'd3730: logsin <= 24'd02056107;
                12'd3731: logsin <= 24'd02056330;
                12'd3732: logsin <= 24'd02056552;
                12'd3733: logsin <= 24'd02056773;
                12'd3734: logsin <= 24'd02056994;
                12'd3735: logsin <= 24'd02057214;
                12'd3736: logsin <= 24'd02057433;
                12'd3737: logsin <= 24'd02057652;
                12'd3738: logsin <= 24'd02057871;
                12'd3739: logsin <= 24'd02058089;
                12'd3740: logsin <= 24'd02058306;
                12'd3741: logsin <= 24'd02058522;
                12'd3742: logsin <= 24'd02058738;
                12'd3743: logsin <= 24'd02058954;
                12'd3744: logsin <= 24'd02059168;
                12'd3745: logsin <= 24'd02059383;
                12'd3746: logsin <= 24'd02059596;
                12'd3747: logsin <= 24'd02059809;
                12'd3748: logsin <= 24'd02060022;
                12'd3749: logsin <= 24'd02060234;
                12'd3750: logsin <= 24'd02060445;
                12'd3751: logsin <= 24'd02060655;
                12'd3752: logsin <= 24'd02060865;
                12'd3753: logsin <= 24'd02061075;
                12'd3754: logsin <= 24'd02061284;
                12'd3755: logsin <= 24'd02061492;
                12'd3756: logsin <= 24'd02061700;
                12'd3757: logsin <= 24'd02061907;
                12'd3758: logsin <= 24'd02062113;
                12'd3759: logsin <= 24'd02062319;
                12'd3760: logsin <= 24'd02062524;
                12'd3761: logsin <= 24'd02062729;
                12'd3762: logsin <= 24'd02062933;
                12'd3763: logsin <= 24'd02063137;
                12'd3764: logsin <= 24'd02063339;
                12'd3765: logsin <= 24'd02063542;
                12'd3766: logsin <= 24'd02063743;
                12'd3767: logsin <= 24'd02063945;
                12'd3768: logsin <= 24'd02064145;
                12'd3769: logsin <= 24'd02064345;
                12'd3770: logsin <= 24'd02064544;
                12'd3771: logsin <= 24'd02064743;
                12'd3772: logsin <= 24'd02064941;
                12'd3773: logsin <= 24'd02065139;
                12'd3774: logsin <= 24'd02065335;
                12'd3775: logsin <= 24'd02065532;
                12'd3776: logsin <= 24'd02065727;
                12'd3777: logsin <= 24'd02065923;
                12'd3778: logsin <= 24'd02066117;
                12'd3779: logsin <= 24'd02066311;
                12'd3780: logsin <= 24'd02066504;
                12'd3781: logsin <= 24'd02066697;
                12'd3782: logsin <= 24'd02066889;
                12'd3783: logsin <= 24'd02067081;
                12'd3784: logsin <= 24'd02067272;
                12'd3785: logsin <= 24'd02067462;
                12'd3786: logsin <= 24'd02067652;
                12'd3787: logsin <= 24'd02067841;
                12'd3788: logsin <= 24'd02068029;
                12'd3789: logsin <= 24'd02068217;
                12'd3790: logsin <= 24'd02068405;
                12'd3791: logsin <= 24'd02068591;
                12'd3792: logsin <= 24'd02068777;
                12'd3793: logsin <= 24'd02068963;
                12'd3794: logsin <= 24'd02069148;
                12'd3795: logsin <= 24'd02069332;
                12'd3796: logsin <= 24'd02069516;
                12'd3797: logsin <= 24'd02069699;
                12'd3798: logsin <= 24'd02069882;
                12'd3799: logsin <= 24'd02070064;
                12'd3800: logsin <= 24'd02070245;
                12'd3801: logsin <= 24'd02070426;
                12'd3802: logsin <= 24'd02070606;
                12'd3803: logsin <= 24'd02070785;
                12'd3804: logsin <= 24'd02070964;
                12'd3805: logsin <= 24'd02071142;
                12'd3806: logsin <= 24'd02071320;
                12'd3807: logsin <= 24'd02071497;
                12'd3808: logsin <= 24'd02071674;
                12'd3809: logsin <= 24'd02071850;
                12'd3810: logsin <= 24'd02072025;
                12'd3811: logsin <= 24'd02072200;
                12'd3812: logsin <= 24'd02072374;
                12'd3813: logsin <= 24'd02072547;
                12'd3814: logsin <= 24'd02072720;
                12'd3815: logsin <= 24'd02072893;
                12'd3816: logsin <= 24'd02073064;
                12'd3817: logsin <= 24'd02073235;
                12'd3818: logsin <= 24'd02073406;
                12'd3819: logsin <= 24'd02073576;
                12'd3820: logsin <= 24'd02073745;
                12'd3821: logsin <= 24'd02073914;
                12'd3822: logsin <= 24'd02074082;
                12'd3823: logsin <= 24'd02074249;
                12'd3824: logsin <= 24'd02074416;
                12'd3825: logsin <= 24'd02074582;
                12'd3826: logsin <= 24'd02074748;
                12'd3827: logsin <= 24'd02074913;
                12'd3828: logsin <= 24'd02075078;
                12'd3829: logsin <= 24'd02075241;
                12'd3830: logsin <= 24'd02075405;
                12'd3831: logsin <= 24'd02075567;
                12'd3832: logsin <= 24'd02075729;
                12'd3833: logsin <= 24'd02075891;
                12'd3834: logsin <= 24'd02076052;
                12'd3835: logsin <= 24'd02076212;
                12'd3836: logsin <= 24'd02076371;
                12'd3837: logsin <= 24'd02076530;
                12'd3838: logsin <= 24'd02076689;
                12'd3839: logsin <= 24'd02076847;
                12'd3840: logsin <= 24'd02077004;
                12'd3841: logsin <= 24'd02077161;
                12'd3842: logsin <= 24'd02077316;
                12'd3843: logsin <= 24'd02077472;
                12'd3844: logsin <= 24'd02077627;
                12'd3845: logsin <= 24'd02077781;
                12'd3846: logsin <= 24'd02077934;
                12'd3847: logsin <= 24'd02078087;
                12'd3848: logsin <= 24'd02078240;
                12'd3849: logsin <= 24'd02078392;
                12'd3850: logsin <= 24'd02078543;
                12'd3851: logsin <= 24'd02078693;
                12'd3852: logsin <= 24'd02078843;
                12'd3853: logsin <= 24'd02078992;
                12'd3854: logsin <= 24'd02079141;
                12'd3855: logsin <= 24'd02079289;
                12'd3856: logsin <= 24'd02079437;
                12'd3857: logsin <= 24'd02079584;
                12'd3858: logsin <= 24'd02079730;
                12'd3859: logsin <= 24'd02079876;
                12'd3860: logsin <= 24'd02080021;
                12'd3861: logsin <= 24'd02080165;
                12'd3862: logsin <= 24'd02080309;
                12'd3863: logsin <= 24'd02080452;
                12'd3864: logsin <= 24'd02080595;
                12'd3865: logsin <= 24'd02080737;
                12'd3866: logsin <= 24'd02080879;
                12'd3867: logsin <= 24'd02081019;
                12'd3868: logsin <= 24'd02081160;
                12'd3869: logsin <= 24'd02081299;
                12'd3870: logsin <= 24'd02081438;
                12'd3871: logsin <= 24'd02081577;
                12'd3872: logsin <= 24'd02081714;
                12'd3873: logsin <= 24'd02081852;
                12'd3874: logsin <= 24'd02081988;
                12'd3875: logsin <= 24'd02082124;
                12'd3876: logsin <= 24'd02082260;
                12'd3877: logsin <= 24'd02082394;
                12'd3878: logsin <= 24'd02082529;
                12'd3879: logsin <= 24'd02082662;
                12'd3880: logsin <= 24'd02082795;
                12'd3881: logsin <= 24'd02082927;
                12'd3882: logsin <= 24'd02083059;
                12'd3883: logsin <= 24'd02083190;
                12'd3884: logsin <= 24'd02083321;
                12'd3885: logsin <= 24'd02083451;
                12'd3886: logsin <= 24'd02083580;
                12'd3887: logsin <= 24'd02083709;
                12'd3888: logsin <= 24'd02083837;
                12'd3889: logsin <= 24'd02083964;
                12'd3890: logsin <= 24'd02084091;
                12'd3891: logsin <= 24'd02084217;
                12'd3892: logsin <= 24'd02084343;
                12'd3893: logsin <= 24'd02084468;
                12'd3894: logsin <= 24'd02084592;
                12'd3895: logsin <= 24'd02084716;
                12'd3896: logsin <= 24'd02084839;
                12'd3897: logsin <= 24'd02084962;
                12'd3898: logsin <= 24'd02085084;
                12'd3899: logsin <= 24'd02085205;
                12'd3900: logsin <= 24'd02085326;
                12'd3901: logsin <= 24'd02085446;
                12'd3902: logsin <= 24'd02085566;
                12'd3903: logsin <= 24'd02085684;
                12'd3904: logsin <= 24'd02085803;
                12'd3905: logsin <= 24'd02085920;
                12'd3906: logsin <= 24'd02086038;
                12'd3907: logsin <= 24'd02086154;
                12'd3908: logsin <= 24'd02086270;
                12'd3909: logsin <= 24'd02086385;
                12'd3910: logsin <= 24'd02086500;
                12'd3911: logsin <= 24'd02086614;
                12'd3912: logsin <= 24'd02086727;
                12'd3913: logsin <= 24'd02086840;
                12'd3914: logsin <= 24'd02086952;
                12'd3915: logsin <= 24'd02087064;
                12'd3916: logsin <= 24'd02087175;
                12'd3917: logsin <= 24'd02087285;
                12'd3918: logsin <= 24'd02087395;
                12'd3919: logsin <= 24'd02087504;
                12'd3920: logsin <= 24'd02087613;
                12'd3921: logsin <= 24'd02087721;
                12'd3922: logsin <= 24'd02087828;
                12'd3923: logsin <= 24'd02087935;
                12'd3924: logsin <= 24'd02088041;
                12'd3925: logsin <= 24'd02088146;
                12'd3926: logsin <= 24'd02088251;
                12'd3927: logsin <= 24'd02088355;
                12'd3928: logsin <= 24'd02088459;
                12'd3929: logsin <= 24'd02088562;
                12'd3930: logsin <= 24'd02088665;
                12'd3931: logsin <= 24'd02088766;
                12'd3932: logsin <= 24'd02088868;
                12'd3933: logsin <= 24'd02088968;
                12'd3934: logsin <= 24'd02089068;
                12'd3935: logsin <= 24'd02089167;
                12'd3936: logsin <= 24'd02089266;
                12'd3937: logsin <= 24'd02089364;
                12'd3938: logsin <= 24'd02089462;
                12'd3939: logsin <= 24'd02089559;
                12'd3940: logsin <= 24'd02089655;
                12'd3941: logsin <= 24'd02089751;
                12'd3942: logsin <= 24'd02089846;
                12'd3943: logsin <= 24'd02089940;
                12'd3944: logsin <= 24'd02090034;
                12'd3945: logsin <= 24'd02090127;
                12'd3946: logsin <= 24'd02090220;
                12'd3947: logsin <= 24'd02090312;
                12'd3948: logsin <= 24'd02090404;
                12'd3949: logsin <= 24'd02090494;
                12'd3950: logsin <= 24'd02090584;
                12'd3951: logsin <= 24'd02090674;
                12'd3952: logsin <= 24'd02090763;
                12'd3953: logsin <= 24'd02090851;
                12'd3954: logsin <= 24'd02090939;
                12'd3955: logsin <= 24'd02091026;
                12'd3956: logsin <= 24'd02091113;
                12'd3957: logsin <= 24'd02091199;
                12'd3958: logsin <= 24'd02091284;
                12'd3959: logsin <= 24'd02091368;
                12'd3960: logsin <= 24'd02091453;
                12'd3961: logsin <= 24'd02091536;
                12'd3962: logsin <= 24'd02091619;
                12'd3963: logsin <= 24'd02091701;
                12'd3964: logsin <= 24'd02091783;
                12'd3965: logsin <= 24'd02091864;
                12'd3966: logsin <= 24'd02091944;
                12'd3967: logsin <= 24'd02092024;
                12'd3968: logsin <= 24'd02092103;
                12'd3969: logsin <= 24'd02092181;
                12'd3970: logsin <= 24'd02092259;
                12'd3971: logsin <= 24'd02092337;
                12'd3972: logsin <= 24'd02092413;
                12'd3973: logsin <= 24'd02092489;
                12'd3974: logsin <= 24'd02092565;
                12'd3975: logsin <= 24'd02092640;
                12'd3976: logsin <= 24'd02092714;
                12'd3977: logsin <= 24'd02092787;
                12'd3978: logsin <= 24'd02092860;
                12'd3979: logsin <= 24'd02092933;
                12'd3980: logsin <= 24'd02093005;
                12'd3981: logsin <= 24'd02093076;
                12'd3982: logsin <= 24'd02093146;
                12'd3983: logsin <= 24'd02093216;
                12'd3984: logsin <= 24'd02093285;
                12'd3985: logsin <= 24'd02093354;
                12'd3986: logsin <= 24'd02093422;
                12'd3987: logsin <= 24'd02093490;
                12'd3988: logsin <= 24'd02093557;
                12'd3989: logsin <= 24'd02093623;
                12'd3990: logsin <= 24'd02093688;
                12'd3991: logsin <= 24'd02093753;
                12'd3992: logsin <= 24'd02093818;
                12'd3993: logsin <= 24'd02093882;
                12'd3994: logsin <= 24'd02093945;
                12'd3995: logsin <= 24'd02094007;
                12'd3996: logsin <= 24'd02094069;
                12'd3997: logsin <= 24'd02094131;
                12'd3998: logsin <= 24'd02094191;
                12'd3999: logsin <= 24'd02094251;
                12'd4000: logsin <= 24'd02094311;
                12'd4001: logsin <= 24'd02094370;
                12'd4002: logsin <= 24'd02094428;
                12'd4003: logsin <= 24'd02094486;
                12'd4004: logsin <= 24'd02094543;
                12'd4005: logsin <= 24'd02094599;
                12'd4006: logsin <= 24'd02094655;
                12'd4007: logsin <= 24'd02094710;
                12'd4008: logsin <= 24'd02094764;
                12'd4009: logsin <= 24'd02094818;
                12'd4010: logsin <= 24'd02094872;
                12'd4011: logsin <= 24'd02094924;
                12'd4012: logsin <= 24'd02094977;
                12'd4013: logsin <= 24'd02095028;
                12'd4014: logsin <= 24'd02095079;
                12'd4015: logsin <= 24'd02095129;
                12'd4016: logsin <= 24'd02095179;
                12'd4017: logsin <= 24'd02095228;
                12'd4018: logsin <= 24'd02095276;
                12'd4019: logsin <= 24'd02095324;
                12'd4020: logsin <= 24'd02095371;
                12'd4021: logsin <= 24'd02095418;
                12'd4022: logsin <= 24'd02095464;
                12'd4023: logsin <= 24'd02095509;
                12'd4024: logsin <= 24'd02095554;
                12'd4025: logsin <= 24'd02095598;
                12'd4026: logsin <= 24'd02095641;
                12'd4027: logsin <= 24'd02095684;
                12'd4028: logsin <= 24'd02095726;
                12'd4029: logsin <= 24'd02095768;
                12'd4030: logsin <= 24'd02095809;
                12'd4031: logsin <= 24'd02095849;
                12'd4032: logsin <= 24'd02095889;
                12'd4033: logsin <= 24'd02095928;
                12'd4034: logsin <= 24'd02095967;
                12'd4035: logsin <= 24'd02096005;
                12'd4036: logsin <= 24'd02096042;
                12'd4037: logsin <= 24'd02096079;
                12'd4038: logsin <= 24'd02096115;
                12'd4039: logsin <= 24'd02096150;
                12'd4040: logsin <= 24'd02096185;
                12'd4041: logsin <= 24'd02096219;
                12'd4042: logsin <= 24'd02096253;
                12'd4043: logsin <= 24'd02096286;
                12'd4044: logsin <= 24'd02096318;
                12'd4045: logsin <= 24'd02096350;
                12'd4046: logsin <= 24'd02096381;
                12'd4047: logsin <= 24'd02096412;
                12'd4048: logsin <= 24'd02096441;
                12'd4049: logsin <= 24'd02096471;
                12'd4050: logsin <= 24'd02096499;
                12'd4051: logsin <= 24'd02096528;
                12'd4052: logsin <= 24'd02096555;
                12'd4053: logsin <= 24'd02096582;
                12'd4054: logsin <= 24'd02096608;
                12'd4055: logsin <= 24'd02096634;
                12'd4056: logsin <= 24'd02096659;
                12'd4057: logsin <= 24'd02096683;
                12'd4058: logsin <= 24'd02096707;
                12'd4059: logsin <= 24'd02096730;
                12'd4060: logsin <= 24'd02096752;
                12'd4061: logsin <= 24'd02096774;
                12'd4062: logsin <= 24'd02096795;
                12'd4063: logsin <= 24'd02096816;
                12'd4064: logsin <= 24'd02096836;
                12'd4065: logsin <= 24'd02096856;
                12'd4066: logsin <= 24'd02096874;
                12'd4067: logsin <= 24'd02096893;
                12'd4068: logsin <= 24'd02096910;
                12'd4069: logsin <= 24'd02096927;
                12'd4070: logsin <= 24'd02096944;
                12'd4071: logsin <= 24'd02096959;
                12'd4072: logsin <= 24'd02096974;
                12'd4073: logsin <= 24'd02096989;
                12'd4074: logsin <= 24'd02097003;
                12'd4075: logsin <= 24'd02097016;
                12'd4076: logsin <= 24'd02097029;
                12'd4077: logsin <= 24'd02097041;
                12'd4078: logsin <= 24'd02097052;
                12'd4079: logsin <= 24'd02097063;
                12'd4080: logsin <= 24'd02097073;
                12'd4081: logsin <= 24'd02097083;
                12'd4082: logsin <= 24'd02097092;
                12'd4083: logsin <= 24'd02097100;
                12'd4084: logsin <= 24'd02097108;
                12'd4085: logsin <= 24'd02097115;
                12'd4086: logsin <= 24'd02097121;
                12'd4087: logsin <= 24'd02097127;
                12'd4088: logsin <= 24'd02097132;
                12'd4089: logsin <= 24'd02097137;
                12'd4090: logsin <= 24'd02097141;
                12'd4091: logsin <= 24'd02097144;
                12'd4092: logsin <= 24'd02097147;
                12'd4093: logsin <= 24'd02097149;
                12'd4094: logsin <= 24'd02097151;
                12'd4095: logsin <= 24'd02097152;
            endcase
        4'b11: //linear512 12/24-bit
            logsin = {3'b000, addr, addr[15:11]};
     
    endcase

endmodule
